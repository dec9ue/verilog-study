

module modexp1 ( e ,n,m, r);
  input[511:0] e,n,m;
  output[511:0] r;

  wire [511:0] m000, r000, 
    m001, r001, m002, r002, m003, r003, m004, r004, m005, r005, m006, r006, m007, r007, m008, r008,
    m009, r009 , m010, r010 , m011, r011 , m012, r012 , m013, r013 , m014, r014 , m015, r015 , m016, r016,
    m017, r017 , m018, r018 , m019, r019 , m020, r020 , m021, r021 , m022, r022 , m023, r023 , m024, r024,
    m025, r025 , m026, r026 , m027, r027 , m028, r028 , m029, r029 , m030, r030 , m031, r031 , m032, r032,
    m033, r033 , m034, r034 , m035, r035 , m036, r036 , m037, r037 , m038, r038 , m039, r039 , m040, r040,
    m041, r041 , m042, r042 , m043, r043 , m044, r044 , m045, r045 , m046, r046 , m047, r047 , m048, r048,
    m049, r049 , m050, r050 , m051, r051 , m052, r052 , m053, r053 , m054, r054 , m055, r055 , m056, r056,
    m057, r057 , m058, r058 , m059, r059 , m060, r060 , m061, r061 , m062, r062 , m063, r063 , m064, r064,
    m065, r065 , m066, r066 , m067, r067 , m068, r068 , m069, r069 , m070, r070 , m071, r071 , m072, r072,
    m073, r073 , m074, r074 , m075, r075 , m076, r076 , m077, r077 , m078, r078 , m079, r079 , m080, r080,
    m081, r081 , m082, r082 , m083, r083 , m084, r084 , m085, r085 , m086, r086 , m087, r087 , m088, r088,
    m089, r089 , m090, r090 , m091, r091 , m092, r092 , m093, r093 , m094, r094 , m095, r095 , m096, r096,
    m097, r097 , m098, r098 , m099, r099 , m100, r100 , m101, r101 , m102, r102 , m103, r103 , m104, r104,
    m105, r105 , m106, r106 , m107, r107 , m108, r108 , m109, r109 , m110, r110 , m111, r111 , m112, r112,
    m113, r113 , m114, r114 , m115, r115 , m116, r116 , m117, r117 , m118, r118 , m119, r119 , m120, r120,
    m121, r121 , m122, r122 , m123, r123 , m124, r124 , m125, r125 , m126, r126 , m127, r127 , m128, r128
    , m129, r129 , m130, r130 , m131, r131 , m132, r132 , m133, r133 , m134, r134 , m135, r135 , m136, r136
    , m137, r137 , m138, r138 , m139, r139 , m140, r140 , m141, r141 , m142, r142 , m143, r143 , m144, r144
    , m145, r145 , m146, r146 , m147, r147 , m148, r148 , m149, r149 , m150, r150 , m151, r151 , m152, r152
    , m153, r153 , m154, r154 , m155, r155 , m156, r156 , m157, r157 , m158, r158 , m159, r159 , m160, r160
    , m161, r161 , m162, r162 , m163, r163 , m164, r164 , m165, r165 , m166, r166 , m167, r167 , m168, r168
    , m169, r169 , m170, r170 , m171, r171 , m172, r172 , m173, r173 , m174, r174 , m175, r175 , m176, r176
    , m177, r177 , m178, r178 , m179, r179 , m180, r180 , m181, r181 , m182, r182 , m183, r183 , m184, r184
    , m185, r185 , m186, r186 , m187, r187 , m188, r188 , m189, r189 , m190, r190 , m191, r191 , m192, r192
    , m193, r193 , m194, r194 , m195, r195 , m196, r196 , m197, r197 , m198, r198 , m199, r199 , m200, r200
    , m201, r201 , m202, r202 , m203, r203 , m204, r204 , m205, r205 , m206, r206 , m207, r207 , m208, r208
    , m209, r209 , m210, r210 , m211, r211 , m212, r212 , m213, r213 , m214, r214 , m215, r215 , m216, r216
    , m217, r217 , m218, r218 , m219, r219 , m220, r220 , m221, r221 , m222, r222 , m223, r223 , m224, r224
    , m225, r225 , m226, r226 , m227, r227 , m228, r228 , m229, r229 , m230, r230 , m231, r231 , m232, r232
    , m233, r233 , m234, r234 , m235, r235 , m236, r236 , m237, r237 , m238, r238 , m239, r239 , m240, r240
    , m241, r241 , m242, r242 , m243, r243 , m244, r244 , m245, r245 , m246, r246 , m247, r247 , m248, r248
    , m249, r249 , m250, r250 , m251, r251 , m252, r252 , m253, r253 , m254, r254 , m255, r255 , m256, r256
    , m257, r257 , m258, r258 , m259, r259 , m260, r260 , m261, r261 , m262, r262 , m263, r263 , m264, r264
    , m265, r265 , m266, r266 , m267, r267 , m268, r268 , m269, r269 , m270, r270 , m271, r271 , m272, r272
    , m273, r273 , m274, r274 , m275, r275 , m276, r276 , m277, r277 , m278, r278 , m279, r279 , m280, r280
    , m281, r281 , m282, r282 , m283, r283 , m284, r284 , m285, r285 , m286, r286 , m287, r287 , m288, r288
    , m289, r289 , m290, r290 , m291, r291 , m292, r292 , m293, r293 , m294, r294 , m295, r295 , m296, r296
    , m297, r297 , m298, r298 , m299, r299 , m300, r300 , m301, r301 , m302, r302 , m303, r303 , m304, r304
    , m305, r305 , m306, r306 , m307, r307 , m308, r308 , m309, r309 , m310, r310 , m311, r311 , m312, r312
    , m313, r313 , m314, r314 , m315, r315 , m316, r316 , m317, r317 , m318, r318 , m319, r319 , m320, r320
    , m321, r321 , m322, r322 , m323, r323 , m324, r324 , m325, r325 , m326, r326 , m327, r327 , m328, r328
    , m329, r329 , m330, r330 , m331, r331 , m332, r332 , m333, r333 , m334, r334 , m335, r335 , m336, r336
    , m337, r337 , m338, r338 , m339, r339 , m340, r340 , m341, r341 , m342, r342 , m343, r343 , m344, r344
    , m345, r345 , m346, r346 , m347, r347 , m348, r348 , m349, r349 , m350, r350 , m351, r351 , m352, r352
    , m353, r353 , m354, r354 , m355, r355 , m356, r356 , m357, r357 , m358, r358 , m359, r359 , m360, r360
    , m361, r361 , m362, r362 , m363, r363 , m364, r364 , m365, r365 , m366, r366 , m367, r367 , m368, r368
    , m369, r369 , m370, r370 , m371, r371 , m372, r372 , m373, r373 , m374, r374 , m375, r375 , m376, r376
    , m377, r377 , m378, r378 , m379, r379 , m380, r380 , m381, r381 , m382, r382 , m383, r383 , m384, r384
    , m385, r385 , m386, r386 , m387, r387 , m388, r388 , m389, r389 , m390, r390 , m391, r391 , m392, r392
    , m393, r393 , m394, r394 , m395, r395 , m396, r396 , m397, r397 , m398, r398 , m399, r399 , m400, r400
    , m401, r401 , m402, r402 , m403, r403 , m404, r404 , m405, r405 , m406, r406 , m407, r407 , m408, r408
    , m409, r409 , m410, r410 , m411, r411 , m412, r412 , m413, r413 , m414, r414 , m415, r415 , m416, r416
    , m417, r417 , m418, r418 , m419, r419 , m420, r420 , m421, r421 , m422, r422 , m423, r423 , m424, r424
    , m425, r425 , m426, r426 , m427, r427 , m428, r428 , m429, r429 , m430, r430 , m431, r431 , m432, r432
    , m433, r433 , m434, r434 , m435, r435 , m436, r436 , m437, r437 , m438, r438 , m439, r439 , m440, r440
    , m441, r441 , m442, r442 , m443, r443 , m444, r444 , m445, r445 , m446, r446 , m447, r447 , m448, r448
    , m449, r449 , m450, r450 , m451, r451 , m452, r452 , m453, r453 , m454, r454 , m455, r455 , m456, r456
    , m457, r457 , m458, r458 , m459, r459 , m460, r460 , m461, r461 , m462, r462 , m463, r463 , m464, r464
    , m465, r465 , m466, r466 , m467, r467 , m468, r468 , m469, r469 , m470, r470 , m471, r471 , m472, r472
    , m473, r473 , m474, r474 , m475, r475 , m476, r476 , m477, r477 , m478, r478 , m479, r479 , m480, r480
    , m481, r481 , m482, r482 , m483, r483 , m484, r484 , m485, r485 , m486, r486 , m487, r487 , m488, r488
    , m489, r489 , m490, r490 , m491, r491 , m492, r492 , m493, r493 , m494, r494 , m495, r495 , m496, r496
    , m497, r497 , m498, r498 , m499, r499 , m500, r500 , m501, r501 , m502, r502 , m503, r503 , m504, r504
    , m505, r505 , m506, r506 , m507, r507 , m508, r508 , m509, r509 , m510, r510 , m511, r511, m512, r512;

  assign m001 = m;
  assign r001 = (1 * (1 + e[0] * (m001 - 1))) % n;

  assign m002 = twice_mod(m001,n); assign r002 = mult_non_zero(r001, e[1],m002) % n;
  assign m003 = twice_mod(m002,n); assign r003 = mult_non_zero(r002, e[2],m003) % n;
  assign m004 = twice_mod(m003,n); assign r004 = mult_non_zero(r003, e[3],m004) % n;
  assign m005 = twice_mod(m004,n); assign r005 = mult_non_zero(r004, e[4],m005) % n;
  assign m006 = twice_mod(m005,n); assign r006 = mult_non_zero(r005, e[5],m006) % n;
  assign m007 = twice_mod(m006,n); assign r007 = mult_non_zero(r006, e[6],m007) % n;
  assign m008 = twice_mod(m007,n); assign r008 = mult_non_zero(r007, e[7],m008) % n;
  assign m009 = twice_mod(m008,n); assign r009 = mult_non_zero(r008, e[8],m009) % n;
  assign m010 = twice_mod(m009,n); assign r010 = mult_non_zero(r009, e[9],m010) % n;
  assign m011 = twice_mod(m010,n); assign r011 = mult_non_zero(r010, e[10],m011) % n;
  assign m012 = twice_mod(m011,n); assign r012 = mult_non_zero(r011, e[11],m012) % n;
  assign m013 = twice_mod(m012,n); assign r013 = mult_non_zero(r012, e[12],m013) % n;
  assign m014 = twice_mod(m013,n); assign r014 = mult_non_zero(r013, e[13],m014) % n;
  assign m015 = twice_mod(m014,n); assign r015 = mult_non_zero(r014, e[14],m015) % n;
  assign m016 = twice_mod(m015,n); assign r016 = mult_non_zero(r015, e[15],m016) % n;
  assign m017 = twice_mod(m016,n); assign r017 = mult_non_zero(r016, e[16],m017) % n;
  assign m018 = twice_mod(m017,n); assign r018 = mult_non_zero(r017, e[17],m018) % n;
  assign m019 = twice_mod(m018,n); assign r019 = mult_non_zero(r018, e[18],m019) % n;
  assign m020 = twice_mod(m019,n); assign r020 = mult_non_zero(r019, e[19],m020) % n;
  assign m021 = twice_mod(m020,n); assign r021 = mult_non_zero(r020, e[20],m021) % n;
  assign m022 = twice_mod(m021,n); assign r022 = mult_non_zero(r021, e[21],m022) % n;
  assign m023 = twice_mod(m022,n); assign r023 = mult_non_zero(r022, e[22],m023) % n;
  assign m024 = twice_mod(m023,n); assign r024 = mult_non_zero(r023, e[23],m024) % n;
  assign m025 = twice_mod(m024,n); assign r025 = mult_non_zero(r024, e[24],m025) % n;
  assign m026 = twice_mod(m025,n); assign r026 = mult_non_zero(r025, e[25],m026) % n;
  assign m027 = twice_mod(m026,n); assign r027 = mult_non_zero(r026, e[26],m027) % n;
  assign m028 = twice_mod(m027,n); assign r028 = mult_non_zero(r027, e[27],m028) % n;
  assign m029 = twice_mod(m028,n); assign r029 = mult_non_zero(r028, e[28],m029) % n;
  assign m030 = twice_mod(m029,n); assign r030 = mult_non_zero(r029, e[29],m030) % n;
  assign m031 = twice_mod(m030,n); assign r031 = mult_non_zero(r030, e[30],m031) % n;
  assign m032 = twice_mod(m031,n); assign r032 = mult_non_zero(r031, e[31],m032) % n;
  assign m033 = twice_mod(m032,n); assign r033 = mult_non_zero(r032, e[32],m033) % n;
  assign m034 = twice_mod(m033,n); assign r034 = mult_non_zero(r033, e[33],m034) % n;
  assign m035 = twice_mod(m034,n); assign r035 = mult_non_zero(r034, e[34],m035) % n;
  assign m036 = twice_mod(m035,n); assign r036 = mult_non_zero(r035, e[35],m036) % n;
  assign m037 = twice_mod(m036,n); assign r037 = mult_non_zero(r036, e[36],m037) % n;
  assign m038 = twice_mod(m037,n); assign r038 = mult_non_zero(r037, e[37],m038) % n;
  assign m039 = twice_mod(m038,n); assign r039 = mult_non_zero(r038, e[38],m039) % n;
  assign m040 = twice_mod(m039,n); assign r040 = mult_non_zero(r039, e[39],m040) % n;
  assign m041 = twice_mod(m040,n); assign r041 = mult_non_zero(r040, e[40],m041) % n;
  assign m042 = twice_mod(m041,n); assign r042 = mult_non_zero(r041, e[41],m042) % n;
  assign m043 = twice_mod(m042,n); assign r043 = mult_non_zero(r042, e[42],m043) % n;
  assign m044 = twice_mod(m043,n); assign r044 = mult_non_zero(r043, e[43],m044) % n;
  assign m045 = twice_mod(m044,n); assign r045 = mult_non_zero(r044, e[44],m045) % n;
  assign m046 = twice_mod(m045,n); assign r046 = mult_non_zero(r045, e[45],m046) % n;
  assign m047 = twice_mod(m046,n); assign r047 = mult_non_zero(r046, e[46],m047) % n;
  assign m048 = twice_mod(m047,n); assign r048 = mult_non_zero(r047, e[47],m048) % n;
  assign m049 = twice_mod(m048,n); assign r049 = mult_non_zero(r048, e[48],m049) % n;
  assign m050 = twice_mod(m049,n); assign r050 = mult_non_zero(r049, e[49],m050) % n;
  assign m051 = twice_mod(m050,n); assign r051 = mult_non_zero(r050, e[50],m051) % n;
  assign m052 = twice_mod(m051,n); assign r052 = mult_non_zero(r051, e[51],m052) % n;
  assign m053 = twice_mod(m052,n); assign r053 = mult_non_zero(r052, e[52],m053) % n;
  assign m054 = twice_mod(m053,n); assign r054 = mult_non_zero(r053, e[53],m054) % n;
  assign m055 = twice_mod(m054,n); assign r055 = mult_non_zero(r054, e[54],m055) % n;
  assign m056 = twice_mod(m055,n); assign r056 = mult_non_zero(r055, e[55],m056) % n;
  assign m057 = twice_mod(m056,n); assign r057 = mult_non_zero(r056, e[56],m057) % n;
  assign m058 = twice_mod(m057,n); assign r058 = mult_non_zero(r057, e[57],m058) % n;
  assign m059 = twice_mod(m058,n); assign r059 = mult_non_zero(r058, e[58],m059) % n;
  assign m060 = twice_mod(m059,n); assign r060 = mult_non_zero(r059, e[59],m060) % n;
  assign m061 = twice_mod(m060,n); assign r061 = mult_non_zero(r060, e[60],m061) % n;
  assign m062 = twice_mod(m061,n); assign r062 = mult_non_zero(r061, e[61],m062) % n;
  assign m063 = twice_mod(m062,n); assign r063 = mult_non_zero(r062, e[62],m063) % n;
  assign m064 = twice_mod(m063,n); assign r064 = mult_non_zero(r063, e[63],m064) % n;
  assign m065 = twice_mod(m064,n); assign r065 = mult_non_zero(r064, e[64],m065) % n;
  assign m066 = twice_mod(m065,n); assign r066 = mult_non_zero(r065, e[65],m066) % n;
  assign m067 = twice_mod(m066,n); assign r067 = mult_non_zero(r066, e[66],m067) % n;
  assign m068 = twice_mod(m067,n); assign r068 = mult_non_zero(r067, e[67],m068) % n;
  assign m069 = twice_mod(m068,n); assign r069 = mult_non_zero(r068, e[68],m069) % n;
  assign m070 = twice_mod(m069,n); assign r070 = mult_non_zero(r069, e[69],m070) % n;
  assign m071 = twice_mod(m070,n); assign r071 = mult_non_zero(r070, e[70],m071) % n;
  assign m072 = twice_mod(m071,n); assign r072 = mult_non_zero(r071, e[71],m072) % n;
  assign m073 = twice_mod(m072,n); assign r073 = mult_non_zero(r072, e[72],m073) % n;
  assign m074 = twice_mod(m073,n); assign r074 = mult_non_zero(r073, e[73],m074) % n;
  assign m075 = twice_mod(m074,n); assign r075 = mult_non_zero(r074, e[74],m075) % n;
  assign m076 = twice_mod(m075,n); assign r076 = mult_non_zero(r075, e[75],m076) % n;
  assign m077 = twice_mod(m076,n); assign r077 = mult_non_zero(r076, e[76],m077) % n;
  assign m078 = twice_mod(m077,n); assign r078 = mult_non_zero(r077, e[77],m078) % n;
  assign m079 = twice_mod(m078,n); assign r079 = mult_non_zero(r078, e[78],m079) % n;
  assign m080 = twice_mod(m079,n); assign r080 = mult_non_zero(r079, e[79],m080) % n;
  assign m081 = twice_mod(m080,n); assign r081 = mult_non_zero(r080, e[80],m081) % n;
  assign m082 = twice_mod(m081,n); assign r082 = mult_non_zero(r081, e[81],m082) % n;
  assign m083 = twice_mod(m082,n); assign r083 = mult_non_zero(r082, e[82],m083) % n;
  assign m084 = twice_mod(m083,n); assign r084 = mult_non_zero(r083, e[83],m084) % n;
  assign m085 = twice_mod(m084,n); assign r085 = mult_non_zero(r084, e[84],m085) % n;
  assign m086 = twice_mod(m085,n); assign r086 = mult_non_zero(r085, e[85],m086) % n;
  assign m087 = twice_mod(m086,n); assign r087 = mult_non_zero(r086, e[86],m087) % n;
  assign m088 = twice_mod(m087,n); assign r088 = mult_non_zero(r087, e[87],m088) % n;
  assign m089 = twice_mod(m088,n); assign r089 = mult_non_zero(r088, e[88],m089) % n;
  assign m090 = twice_mod(m089,n); assign r090 = mult_non_zero(r089, e[89],m090) % n;
  assign m091 = twice_mod(m090,n); assign r091 = mult_non_zero(r090, e[90],m091) % n;
  assign m092 = twice_mod(m091,n); assign r092 = mult_non_zero(r091, e[91],m092) % n;
  assign m093 = twice_mod(m092,n); assign r093 = mult_non_zero(r092, e[92],m093) % n;
  assign m094 = twice_mod(m093,n); assign r094 = mult_non_zero(r093, e[93],m094) % n;
  assign m095 = twice_mod(m094,n); assign r095 = mult_non_zero(r094, e[94],m095) % n;
  assign m096 = twice_mod(m095,n); assign r096 = mult_non_zero(r095, e[95],m096) % n;
  assign m097 = twice_mod(m096,n); assign r097 = mult_non_zero(r096, e[96],m097) % n;
  assign m098 = twice_mod(m097,n); assign r098 = mult_non_zero(r097, e[97],m098) % n;
  assign m099 = twice_mod(m098,n); assign r099 = mult_non_zero(r098, e[98],m099) % n;
  assign m100 = twice_mod(m099,n); assign r100 = mult_non_zero(r099, e[99],m100) % n;
  assign m101 = twice_mod(m100,n); assign r101 = mult_non_zero(r100, e[100],m101) % n;
  assign m102 = twice_mod(m101,n); assign r102 = mult_non_zero(r101, e[101],m102) % n;
  assign m103 = twice_mod(m102,n); assign r103 = mult_non_zero(r102, e[102],m103) % n;
  assign m104 = twice_mod(m103,n); assign r104 = mult_non_zero(r103, e[103],m104) % n;
  assign m105 = twice_mod(m104,n); assign r105 = mult_non_zero(r104, e[104],m105) % n;
  assign m106 = twice_mod(m105,n); assign r106 = mult_non_zero(r105, e[105],m106) % n;
  assign m107 = twice_mod(m106,n); assign r107 = mult_non_zero(r106, e[106],m107) % n;
  assign m108 = twice_mod(m107,n); assign r108 = mult_non_zero(r107, e[107],m108) % n;
  assign m109 = twice_mod(m108,n); assign r109 = mult_non_zero(r108, e[108],m109) % n;
  assign m110 = twice_mod(m109,n); assign r110 = mult_non_zero(r109, e[109],m110) % n;
  assign m111 = twice_mod(m110,n); assign r111 = mult_non_zero(r110, e[110],m111) % n;
  assign m112 = twice_mod(m111,n); assign r112 = mult_non_zero(r111, e[111],m112) % n;
  assign m113 = twice_mod(m112,n); assign r113 = mult_non_zero(r112, e[112],m113) % n;
  assign m114 = twice_mod(m113,n); assign r114 = mult_non_zero(r113, e[113],m114) % n;
  assign m115 = twice_mod(m114,n); assign r115 = mult_non_zero(r114, e[114],m115) % n;
  assign m116 = twice_mod(m115,n); assign r116 = mult_non_zero(r115, e[115],m116) % n;
  assign m117 = twice_mod(m116,n); assign r117 = mult_non_zero(r116, e[116],m117) % n;
  assign m118 = twice_mod(m117,n); assign r118 = mult_non_zero(r117, e[117],m118) % n;
  assign m119 = twice_mod(m118,n); assign r119 = mult_non_zero(r118, e[118],m119) % n;
  assign m120 = twice_mod(m119,n); assign r120 = mult_non_zero(r119, e[119],m120) % n;
  assign m121 = twice_mod(m120,n); assign r121 = mult_non_zero(r120, e[120],m121) % n;
  assign m122 = twice_mod(m121,n); assign r122 = mult_non_zero(r121, e[121],m122) % n;
  assign m123 = twice_mod(m122,n); assign r123 = mult_non_zero(r122, e[122],m123) % n;
  assign m124 = twice_mod(m123,n); assign r124 = mult_non_zero(r123, e[123],m124) % n;
  assign m125 = twice_mod(m124,n); assign r125 = mult_non_zero(r124, e[124],m125) % n;
  assign m126 = twice_mod(m125,n); assign r126 = mult_non_zero(r125, e[125],m126) % n;
  assign m127 = twice_mod(m126,n); assign r127 = mult_non_zero(r126, e[126],m127) % n;
  assign m128 = twice_mod(m127,n); assign r128 = mult_non_zero(r127, e[127],m128) % n;
  assign m129 = twice_mod(m128,n); assign r129 = mult_non_zero(r128, e[128],m129) % n;
  assign m130 = twice_mod(m129,n); assign r130 = mult_non_zero(r129, e[129],m130) % n;
  assign m131 = twice_mod(m130,n); assign r131 = mult_non_zero(r130, e[130],m131) % n;
  assign m132 = twice_mod(m131,n); assign r132 = mult_non_zero(r131, e[131],m132) % n;
  assign m133 = twice_mod(m132,n); assign r133 = mult_non_zero(r132, e[132],m133) % n;
  assign m134 = twice_mod(m133,n); assign r134 = mult_non_zero(r133, e[133],m134) % n;
  assign m135 = twice_mod(m134,n); assign r135 = mult_non_zero(r134, e[134],m135) % n;
  assign m136 = twice_mod(m135,n); assign r136 = mult_non_zero(r135, e[135],m136) % n;
  assign m137 = twice_mod(m136,n); assign r137 = mult_non_zero(r136, e[136],m137) % n;
  assign m138 = twice_mod(m137,n); assign r138 = mult_non_zero(r137, e[137],m138) % n;
  assign m139 = twice_mod(m138,n); assign r139 = mult_non_zero(r138, e[138],m139) % n;
  assign m140 = twice_mod(m139,n); assign r140 = mult_non_zero(r139, e[139],m140) % n;
  assign m141 = twice_mod(m140,n); assign r141 = mult_non_zero(r140, e[140],m141) % n;
  assign m142 = twice_mod(m141,n); assign r142 = mult_non_zero(r141, e[141],m142) % n;
  assign m143 = twice_mod(m142,n); assign r143 = mult_non_zero(r142, e[142],m143) % n;
  assign m144 = twice_mod(m143,n); assign r144 = mult_non_zero(r143, e[143],m144) % n;
  assign m145 = twice_mod(m144,n); assign r145 = mult_non_zero(r144, e[144],m145) % n;
  assign m146 = twice_mod(m145,n); assign r146 = mult_non_zero(r145, e[145],m146) % n;
  assign m147 = twice_mod(m146,n); assign r147 = mult_non_zero(r146, e[146],m147) % n;
  assign m148 = twice_mod(m147,n); assign r148 = mult_non_zero(r147, e[147],m148) % n;
  assign m149 = twice_mod(m148,n); assign r149 = mult_non_zero(r148, e[148],m149) % n;
  assign m150 = twice_mod(m149,n); assign r150 = mult_non_zero(r149, e[149],m150) % n;
  assign m151 = twice_mod(m150,n); assign r151 = mult_non_zero(r150, e[150],m151) % n;
  assign m152 = twice_mod(m151,n); assign r152 = mult_non_zero(r151, e[151],m152) % n;
  assign m153 = twice_mod(m152,n); assign r153 = mult_non_zero(r152, e[152],m153) % n;
  assign m154 = twice_mod(m153,n); assign r154 = mult_non_zero(r153, e[153],m154) % n;
  assign m155 = twice_mod(m154,n); assign r155 = mult_non_zero(r154, e[154],m155) % n;
  assign m156 = twice_mod(m155,n); assign r156 = mult_non_zero(r155, e[155],m156) % n;
  assign m157 = twice_mod(m156,n); assign r157 = mult_non_zero(r156, e[156],m157) % n;
  assign m158 = twice_mod(m157,n); assign r158 = mult_non_zero(r157, e[157],m158) % n;
  assign m159 = twice_mod(m158,n); assign r159 = mult_non_zero(r158, e[158],m159) % n;
  assign m160 = twice_mod(m159,n); assign r160 = mult_non_zero(r159, e[159],m160) % n;
  assign m161 = twice_mod(m160,n); assign r161 = mult_non_zero(r160, e[160],m161) % n;
  assign m162 = twice_mod(m161,n); assign r162 = mult_non_zero(r161, e[161],m162) % n;
  assign m163 = twice_mod(m162,n); assign r163 = mult_non_zero(r162, e[162],m163) % n;
  assign m164 = twice_mod(m163,n); assign r164 = mult_non_zero(r163, e[163],m164) % n;
  assign m165 = twice_mod(m164,n); assign r165 = mult_non_zero(r164, e[164],m165) % n;
  assign m166 = twice_mod(m165,n); assign r166 = mult_non_zero(r165, e[165],m166) % n;
  assign m167 = twice_mod(m166,n); assign r167 = mult_non_zero(r166, e[166],m167) % n;
  assign m168 = twice_mod(m167,n); assign r168 = mult_non_zero(r167, e[167],m168) % n;
  assign m169 = twice_mod(m168,n); assign r169 = mult_non_zero(r168, e[168],m169) % n;
  assign m170 = twice_mod(m169,n); assign r170 = mult_non_zero(r169, e[169],m170) % n;
  assign m171 = twice_mod(m170,n); assign r171 = mult_non_zero(r170, e[170],m171) % n;
  assign m172 = twice_mod(m171,n); assign r172 = mult_non_zero(r171, e[171],m172) % n;
  assign m173 = twice_mod(m172,n); assign r173 = mult_non_zero(r172, e[172],m173) % n;
  assign m174 = twice_mod(m173,n); assign r174 = mult_non_zero(r173, e[173],m174) % n;
  assign m175 = twice_mod(m174,n); assign r175 = mult_non_zero(r174, e[174],m175) % n;
  assign m176 = twice_mod(m175,n); assign r176 = mult_non_zero(r175, e[175],m176) % n;
  assign m177 = twice_mod(m176,n); assign r177 = mult_non_zero(r176, e[176],m177) % n;
  assign m178 = twice_mod(m177,n); assign r178 = mult_non_zero(r177, e[177],m178) % n;
  assign m179 = twice_mod(m178,n); assign r179 = mult_non_zero(r178, e[178],m179) % n;
  assign m180 = twice_mod(m179,n); assign r180 = mult_non_zero(r179, e[179],m180) % n;
  assign m181 = twice_mod(m180,n); assign r181 = mult_non_zero(r180, e[180],m181) % n;
  assign m182 = twice_mod(m181,n); assign r182 = mult_non_zero(r181, e[181],m182) % n;
  assign m183 = twice_mod(m182,n); assign r183 = mult_non_zero(r182, e[182],m183) % n;
  assign m184 = twice_mod(m183,n); assign r184 = mult_non_zero(r183, e[183],m184) % n;
  assign m185 = twice_mod(m184,n); assign r185 = mult_non_zero(r184, e[184],m185) % n;
  assign m186 = twice_mod(m185,n); assign r186 = mult_non_zero(r185, e[185],m186) % n;
  assign m187 = twice_mod(m186,n); assign r187 = mult_non_zero(r186, e[186],m187) % n;
  assign m188 = twice_mod(m187,n); assign r188 = mult_non_zero(r187, e[187],m188) % n;
  assign m189 = twice_mod(m188,n); assign r189 = mult_non_zero(r188, e[188],m189) % n;
  assign m190 = twice_mod(m189,n); assign r190 = mult_non_zero(r189, e[189],m190) % n;
  assign m191 = twice_mod(m190,n); assign r191 = mult_non_zero(r190, e[190],m191) % n;
  assign m192 = twice_mod(m191,n); assign r192 = mult_non_zero(r191, e[191],m192) % n;
  assign m193 = twice_mod(m192,n); assign r193 = mult_non_zero(r192, e[192],m193) % n;
  assign m194 = twice_mod(m193,n); assign r194 = mult_non_zero(r193, e[193],m194) % n;
  assign m195 = twice_mod(m194,n); assign r195 = mult_non_zero(r194, e[194],m195) % n;
  assign m196 = twice_mod(m195,n); assign r196 = mult_non_zero(r195, e[195],m196) % n;
  assign m197 = twice_mod(m196,n); assign r197 = mult_non_zero(r196, e[196],m197) % n;
  assign m198 = twice_mod(m197,n); assign r198 = mult_non_zero(r197, e[197],m198) % n;
  assign m199 = twice_mod(m198,n); assign r199 = mult_non_zero(r198, e[198],m199) % n;
  assign m200 = twice_mod(m199,n); assign r200 = mult_non_zero(r199, e[199],m200) % n;
  assign m201 = twice_mod(m200,n); assign r201 = mult_non_zero(r200, e[200],m201) % n;
  assign m202 = twice_mod(m201,n); assign r202 = mult_non_zero(r201, e[201],m202) % n;
  assign m203 = twice_mod(m202,n); assign r203 = mult_non_zero(r202, e[202],m203) % n;
  assign m204 = twice_mod(m203,n); assign r204 = mult_non_zero(r203, e[203],m204) % n;
  assign m205 = twice_mod(m204,n); assign r205 = mult_non_zero(r204, e[204],m205) % n;
  assign m206 = twice_mod(m205,n); assign r206 = mult_non_zero(r205, e[205],m206) % n;
  assign m207 = twice_mod(m206,n); assign r207 = mult_non_zero(r206, e[206],m207) % n;
  assign m208 = twice_mod(m207,n); assign r208 = mult_non_zero(r207, e[207],m208) % n;
  assign m209 = twice_mod(m208,n); assign r209 = mult_non_zero(r208, e[208],m209) % n;
  assign m210 = twice_mod(m209,n); assign r210 = mult_non_zero(r209, e[209],m210) % n;
  assign m211 = twice_mod(m210,n); assign r211 = mult_non_zero(r210, e[210],m211) % n;
  assign m212 = twice_mod(m211,n); assign r212 = mult_non_zero(r211, e[211],m212) % n;
  assign m213 = twice_mod(m212,n); assign r213 = mult_non_zero(r212, e[212],m213) % n;
  assign m214 = twice_mod(m213,n); assign r214 = mult_non_zero(r213, e[213],m214) % n;
  assign m215 = twice_mod(m214,n); assign r215 = mult_non_zero(r214, e[214],m215) % n;
  assign m216 = twice_mod(m215,n); assign r216 = mult_non_zero(r215, e[215],m216) % n;
  assign m217 = twice_mod(m216,n); assign r217 = mult_non_zero(r216, e[216],m217) % n;
  assign m218 = twice_mod(m217,n); assign r218 = mult_non_zero(r217, e[217],m218) % n;
  assign m219 = twice_mod(m218,n); assign r219 = mult_non_zero(r218, e[218],m219) % n;
  assign m220 = twice_mod(m219,n); assign r220 = mult_non_zero(r219, e[219],m220) % n;
  assign m221 = twice_mod(m220,n); assign r221 = mult_non_zero(r220, e[220],m221) % n;
  assign m222 = twice_mod(m221,n); assign r222 = mult_non_zero(r221, e[221],m222) % n;
  assign m223 = twice_mod(m222,n); assign r223 = mult_non_zero(r222, e[222],m223) % n;
  assign m224 = twice_mod(m223,n); assign r224 = mult_non_zero(r223, e[223],m224) % n;
  assign m225 = twice_mod(m224,n); assign r225 = mult_non_zero(r224, e[224],m225) % n;
  assign m226 = twice_mod(m225,n); assign r226 = mult_non_zero(r225, e[225],m226) % n;
  assign m227 = twice_mod(m226,n); assign r227 = mult_non_zero(r226, e[226],m227) % n;
  assign m228 = twice_mod(m227,n); assign r228 = mult_non_zero(r227, e[227],m228) % n;
  assign m229 = twice_mod(m228,n); assign r229 = mult_non_zero(r228, e[228],m229) % n;
  assign m230 = twice_mod(m229,n); assign r230 = mult_non_zero(r229, e[229],m230) % n;
  assign m231 = twice_mod(m230,n); assign r231 = mult_non_zero(r230, e[230],m231) % n;
  assign m232 = twice_mod(m231,n); assign r232 = mult_non_zero(r231, e[231],m232) % n;
  assign m233 = twice_mod(m232,n); assign r233 = mult_non_zero(r232, e[232],m233) % n;
  assign m234 = twice_mod(m233,n); assign r234 = mult_non_zero(r233, e[233],m234) % n;
  assign m235 = twice_mod(m234,n); assign r235 = mult_non_zero(r234, e[234],m235) % n;
  assign m236 = twice_mod(m235,n); assign r236 = mult_non_zero(r235, e[235],m236) % n;
  assign m237 = twice_mod(m236,n); assign r237 = mult_non_zero(r236, e[236],m237) % n;
  assign m238 = twice_mod(m237,n); assign r238 = mult_non_zero(r237, e[237],m238) % n;
  assign m239 = twice_mod(m238,n); assign r239 = mult_non_zero(r238, e[238],m239) % n;
  assign m240 = twice_mod(m239,n); assign r240 = mult_non_zero(r239, e[239],m240) % n;
  assign m241 = twice_mod(m240,n); assign r241 = mult_non_zero(r240, e[240],m241) % n;
  assign m242 = twice_mod(m241,n); assign r242 = mult_non_zero(r241, e[241],m242) % n;
  assign m243 = twice_mod(m242,n); assign r243 = mult_non_zero(r242, e[242],m243) % n;
  assign m244 = twice_mod(m243,n); assign r244 = mult_non_zero(r243, e[243],m244) % n;
  assign m245 = twice_mod(m244,n); assign r245 = mult_non_zero(r244, e[244],m245) % n;
  assign m246 = twice_mod(m245,n); assign r246 = mult_non_zero(r245, e[245],m246) % n;
  assign m247 = twice_mod(m246,n); assign r247 = mult_non_zero(r246, e[246],m247) % n;
  assign m248 = twice_mod(m247,n); assign r248 = mult_non_zero(r247, e[247],m248) % n;
  assign m249 = twice_mod(m248,n); assign r249 = mult_non_zero(r248, e[248],m249) % n;
  assign m250 = twice_mod(m249,n); assign r250 = mult_non_zero(r249, e[249],m250) % n;
  assign m251 = twice_mod(m250,n); assign r251 = mult_non_zero(r250, e[250],m251) % n;
  assign m252 = twice_mod(m251,n); assign r252 = mult_non_zero(r251, e[251],m252) % n;
  assign m253 = twice_mod(m252,n); assign r253 = mult_non_zero(r252, e[252],m253) % n;
  assign m254 = twice_mod(m253,n); assign r254 = mult_non_zero(r253, e[253],m254) % n;
  assign m255 = twice_mod(m254,n); assign r255 = mult_non_zero(r254, e[254],m255) % n;
  assign m256 = twice_mod(m255,n); assign r256 = mult_non_zero(r255, e[255],m256) % n;
  assign m257 = twice_mod(m256,n); assign r257 = mult_non_zero(r256, e[256],m257) % n;
  assign m258 = twice_mod(m257,n); assign r258 = mult_non_zero(r257, e[257],m258) % n;
  assign m259 = twice_mod(m258,n); assign r259 = mult_non_zero(r258, e[258],m259) % n;
  assign m260 = twice_mod(m259,n); assign r260 = mult_non_zero(r259, e[259],m260) % n;
  assign m261 = twice_mod(m260,n); assign r261 = mult_non_zero(r260, e[260],m261) % n;
  assign m262 = twice_mod(m261,n); assign r262 = mult_non_zero(r261, e[261],m262) % n;
  assign m263 = twice_mod(m262,n); assign r263 = mult_non_zero(r262, e[262],m263) % n;
  assign m264 = twice_mod(m263,n); assign r264 = mult_non_zero(r263, e[263],m264) % n;
  assign m265 = twice_mod(m264,n); assign r265 = mult_non_zero(r264, e[264],m265) % n;
  assign m266 = twice_mod(m265,n); assign r266 = mult_non_zero(r265, e[265],m266) % n;
  assign m267 = twice_mod(m266,n); assign r267 = mult_non_zero(r266, e[266],m267) % n;
  assign m268 = twice_mod(m267,n); assign r268 = mult_non_zero(r267, e[267],m268) % n;
  assign m269 = twice_mod(m268,n); assign r269 = mult_non_zero(r268, e[268],m269) % n;
  assign m270 = twice_mod(m269,n); assign r270 = mult_non_zero(r269, e[269],m270) % n;
  assign m271 = twice_mod(m270,n); assign r271 = mult_non_zero(r270, e[270],m271) % n;
  assign m272 = twice_mod(m271,n); assign r272 = mult_non_zero(r271, e[271],m272) % n;
  assign m273 = twice_mod(m272,n); assign r273 = mult_non_zero(r272, e[272],m273) % n;
  assign m274 = twice_mod(m273,n); assign r274 = mult_non_zero(r273, e[273],m274) % n;
  assign m275 = twice_mod(m274,n); assign r275 = mult_non_zero(r274, e[274],m275) % n;
  assign m276 = twice_mod(m275,n); assign r276 = mult_non_zero(r275, e[275],m276) % n;
  assign m277 = twice_mod(m276,n); assign r277 = mult_non_zero(r276, e[276],m277) % n;
  assign m278 = twice_mod(m277,n); assign r278 = mult_non_zero(r277, e[277],m278) % n;
  assign m279 = twice_mod(m278,n); assign r279 = mult_non_zero(r278, e[278],m279) % n;
  assign m280 = twice_mod(m279,n); assign r280 = mult_non_zero(r279, e[279],m280) % n;
  assign m281 = twice_mod(m280,n); assign r281 = mult_non_zero(r280, e[280],m281) % n;
  assign m282 = twice_mod(m281,n); assign r282 = mult_non_zero(r281, e[281],m282) % n;
  assign m283 = twice_mod(m282,n); assign r283 = mult_non_zero(r282, e[282],m283) % n;
  assign m284 = twice_mod(m283,n); assign r284 = mult_non_zero(r283, e[283],m284) % n;
  assign m285 = twice_mod(m284,n); assign r285 = mult_non_zero(r284, e[284],m285) % n;
  assign m286 = twice_mod(m285,n); assign r286 = mult_non_zero(r285, e[285],m286) % n;
  assign m287 = twice_mod(m286,n); assign r287 = mult_non_zero(r286, e[286],m287) % n;
  assign m288 = twice_mod(m287,n); assign r288 = mult_non_zero(r287, e[287],m288) % n;
  assign m289 = twice_mod(m288,n); assign r289 = mult_non_zero(r288, e[288],m289) % n;
  assign m290 = twice_mod(m289,n); assign r290 = mult_non_zero(r289, e[289],m290) % n;
  assign m291 = twice_mod(m290,n); assign r291 = mult_non_zero(r290, e[290],m291) % n;
  assign m292 = twice_mod(m291,n); assign r292 = mult_non_zero(r291, e[291],m292) % n;
  assign m293 = twice_mod(m292,n); assign r293 = mult_non_zero(r292, e[292],m293) % n;
  assign m294 = twice_mod(m293,n); assign r294 = mult_non_zero(r293, e[293],m294) % n;
  assign m295 = twice_mod(m294,n); assign r295 = mult_non_zero(r294, e[294],m295) % n;
  assign m296 = twice_mod(m295,n); assign r296 = mult_non_zero(r295, e[295],m296) % n;
  assign m297 = twice_mod(m296,n); assign r297 = mult_non_zero(r296, e[296],m297) % n;
  assign m298 = twice_mod(m297,n); assign r298 = mult_non_zero(r297, e[297],m298) % n;
  assign m299 = twice_mod(m298,n); assign r299 = mult_non_zero(r298, e[298],m299) % n;
  assign m300 = twice_mod(m299,n); assign r300 = mult_non_zero(r299, e[299],m300) % n;
  assign m301 = twice_mod(m300,n); assign r301 = mult_non_zero(r300, e[300],m301) % n;
  assign m302 = twice_mod(m301,n); assign r302 = mult_non_zero(r301, e[301],m302) % n;
  assign m303 = twice_mod(m302,n); assign r303 = mult_non_zero(r302, e[302],m303) % n;
  assign m304 = twice_mod(m303,n); assign r304 = mult_non_zero(r303, e[303],m304) % n;
  assign m305 = twice_mod(m304,n); assign r305 = mult_non_zero(r304, e[304],m305) % n;
  assign m306 = twice_mod(m305,n); assign r306 = mult_non_zero(r305, e[305],m306) % n;
  assign m307 = twice_mod(m306,n); assign r307 = mult_non_zero(r306, e[306],m307) % n;
  assign m308 = twice_mod(m307,n); assign r308 = mult_non_zero(r307, e[307],m308) % n;
  assign m309 = twice_mod(m308,n); assign r309 = mult_non_zero(r308, e[308],m309) % n;
  assign m310 = twice_mod(m309,n); assign r310 = mult_non_zero(r309, e[309],m310) % n;
  assign m311 = twice_mod(m310,n); assign r311 = mult_non_zero(r310, e[310],m311) % n;
  assign m312 = twice_mod(m311,n); assign r312 = mult_non_zero(r311, e[311],m312) % n;
  assign m313 = twice_mod(m312,n); assign r313 = mult_non_zero(r312, e[312],m313) % n;
  assign m314 = twice_mod(m313,n); assign r314 = mult_non_zero(r313, e[313],m314) % n;
  assign m315 = twice_mod(m314,n); assign r315 = mult_non_zero(r314, e[314],m315) % n;
  assign m316 = twice_mod(m315,n); assign r316 = mult_non_zero(r315, e[315],m316) % n;
  assign m317 = twice_mod(m316,n); assign r317 = mult_non_zero(r316, e[316],m317) % n;
  assign m318 = twice_mod(m317,n); assign r318 = mult_non_zero(r317, e[317],m318) % n;
  assign m319 = twice_mod(m318,n); assign r319 = mult_non_zero(r318, e[318],m319) % n;
  assign m320 = twice_mod(m319,n); assign r320 = mult_non_zero(r319, e[319],m320) % n;
  assign m321 = twice_mod(m320,n); assign r321 = mult_non_zero(r320, e[320],m321) % n;
  assign m322 = twice_mod(m321,n); assign r322 = mult_non_zero(r321, e[321],m322) % n;
  assign m323 = twice_mod(m322,n); assign r323 = mult_non_zero(r322, e[322],m323) % n;
  assign m324 = twice_mod(m323,n); assign r324 = mult_non_zero(r323, e[323],m324) % n;
  assign m325 = twice_mod(m324,n); assign r325 = mult_non_zero(r324, e[324],m325) % n;
  assign m326 = twice_mod(m325,n); assign r326 = mult_non_zero(r325, e[325],m326) % n;
  assign m327 = twice_mod(m326,n); assign r327 = mult_non_zero(r326, e[326],m327) % n;
  assign m328 = twice_mod(m327,n); assign r328 = mult_non_zero(r327, e[327],m328) % n;
  assign m329 = twice_mod(m328,n); assign r329 = mult_non_zero(r328, e[328],m329) % n;
  assign m330 = twice_mod(m329,n); assign r330 = mult_non_zero(r329, e[329],m330) % n;
  assign m331 = twice_mod(m330,n); assign r331 = mult_non_zero(r330, e[330],m331) % n;
  assign m332 = twice_mod(m331,n); assign r332 = mult_non_zero(r331, e[331],m332) % n;
  assign m333 = twice_mod(m332,n); assign r333 = mult_non_zero(r332, e[332],m333) % n;
  assign m334 = twice_mod(m333,n); assign r334 = mult_non_zero(r333, e[333],m334) % n;
  assign m335 = twice_mod(m334,n); assign r335 = mult_non_zero(r334, e[334],m335) % n;
  assign m336 = twice_mod(m335,n); assign r336 = mult_non_zero(r335, e[335],m336) % n;
  assign m337 = twice_mod(m336,n); assign r337 = mult_non_zero(r336, e[336],m337) % n;
  assign m338 = twice_mod(m337,n); assign r338 = mult_non_zero(r337, e[337],m338) % n;
  assign m339 = twice_mod(m338,n); assign r339 = mult_non_zero(r338, e[338],m339) % n;
  assign m340 = twice_mod(m339,n); assign r340 = mult_non_zero(r339, e[339],m340) % n;
  assign m341 = twice_mod(m340,n); assign r341 = mult_non_zero(r340, e[340],m341) % n;
  assign m342 = twice_mod(m341,n); assign r342 = mult_non_zero(r341, e[341],m342) % n;
  assign m343 = twice_mod(m342,n); assign r343 = mult_non_zero(r342, e[342],m343) % n;
  assign m344 = twice_mod(m343,n); assign r344 = mult_non_zero(r343, e[343],m344) % n;
  assign m345 = twice_mod(m344,n); assign r345 = mult_non_zero(r344, e[344],m345) % n;
  assign m346 = twice_mod(m345,n); assign r346 = mult_non_zero(r345, e[345],m346) % n;
  assign m347 = twice_mod(m346,n); assign r347 = mult_non_zero(r346, e[346],m347) % n;
  assign m348 = twice_mod(m347,n); assign r348 = mult_non_zero(r347, e[347],m348) % n;
  assign m349 = twice_mod(m348,n); assign r349 = mult_non_zero(r348, e[348],m349) % n;
  assign m350 = twice_mod(m349,n); assign r350 = mult_non_zero(r349, e[349],m350) % n;
  assign m351 = twice_mod(m350,n); assign r351 = mult_non_zero(r350, e[350],m351) % n;
  assign m352 = twice_mod(m351,n); assign r352 = mult_non_zero(r351, e[351],m352) % n;
  assign m353 = twice_mod(m352,n); assign r353 = mult_non_zero(r352, e[352],m353) % n;
  assign m354 = twice_mod(m353,n); assign r354 = mult_non_zero(r353, e[353],m354) % n;
  assign m355 = twice_mod(m354,n); assign r355 = mult_non_zero(r354, e[354],m355) % n;
  assign m356 = twice_mod(m355,n); assign r356 = mult_non_zero(r355, e[355],m356) % n;
  assign m357 = twice_mod(m356,n); assign r357 = mult_non_zero(r356, e[356],m357) % n;
  assign m358 = twice_mod(m357,n); assign r358 = mult_non_zero(r357, e[357],m358) % n;
  assign m359 = twice_mod(m358,n); assign r359 = mult_non_zero(r358, e[358],m359) % n;
  assign m360 = twice_mod(m359,n); assign r360 = mult_non_zero(r359, e[359],m360) % n;
  assign m361 = twice_mod(m360,n); assign r361 = mult_non_zero(r360, e[360],m361) % n;
  assign m362 = twice_mod(m361,n); assign r362 = mult_non_zero(r361, e[361],m362) % n;
  assign m363 = twice_mod(m362,n); assign r363 = mult_non_zero(r362, e[362],m363) % n;
  assign m364 = twice_mod(m363,n); assign r364 = mult_non_zero(r363, e[363],m364) % n;
  assign m365 = twice_mod(m364,n); assign r365 = mult_non_zero(r364, e[364],m365) % n;
  assign m366 = twice_mod(m365,n); assign r366 = mult_non_zero(r365, e[365],m366) % n;
  assign m367 = twice_mod(m366,n); assign r367 = mult_non_zero(r366, e[366],m367) % n;
  assign m368 = twice_mod(m367,n); assign r368 = mult_non_zero(r367, e[367],m368) % n;
  assign m369 = twice_mod(m368,n); assign r369 = mult_non_zero(r368, e[368],m369) % n;
  assign m370 = twice_mod(m369,n); assign r370 = mult_non_zero(r369, e[369],m370) % n;
  assign m371 = twice_mod(m370,n); assign r371 = mult_non_zero(r370, e[370],m371) % n;
  assign m372 = twice_mod(m371,n); assign r372 = mult_non_zero(r371, e[371],m372) % n;
  assign m373 = twice_mod(m372,n); assign r373 = mult_non_zero(r372, e[372],m373) % n;
  assign m374 = twice_mod(m373,n); assign r374 = mult_non_zero(r373, e[373],m374) % n;
  assign m375 = twice_mod(m374,n); assign r375 = mult_non_zero(r374, e[374],m375) % n;
  assign m376 = twice_mod(m375,n); assign r376 = mult_non_zero(r375, e[375],m376) % n;
  assign m377 = twice_mod(m376,n); assign r377 = mult_non_zero(r376, e[376],m377) % n;
  assign m378 = twice_mod(m377,n); assign r378 = mult_non_zero(r377, e[377],m378) % n;
  assign m379 = twice_mod(m378,n); assign r379 = mult_non_zero(r378, e[378],m379) % n;
  assign m380 = twice_mod(m379,n); assign r380 = mult_non_zero(r379, e[379],m380) % n;
  assign m381 = twice_mod(m380,n); assign r381 = mult_non_zero(r380, e[380],m381) % n;
  assign m382 = twice_mod(m381,n); assign r382 = mult_non_zero(r381, e[381],m382) % n;
  assign m383 = twice_mod(m382,n); assign r383 = mult_non_zero(r382, e[382],m383) % n;
  assign m384 = twice_mod(m383,n); assign r384 = mult_non_zero(r383, e[383],m384) % n;
  assign m385 = twice_mod(m384,n); assign r385 = mult_non_zero(r384, e[384],m385) % n;
  assign m386 = twice_mod(m385,n); assign r386 = mult_non_zero(r385, e[385],m386) % n;
  assign m387 = twice_mod(m386,n); assign r387 = mult_non_zero(r386, e[386],m387) % n;
  assign m388 = twice_mod(m387,n); assign r388 = mult_non_zero(r387, e[387],m388) % n;
  assign m389 = twice_mod(m388,n); assign r389 = mult_non_zero(r388, e[388],m389) % n;
  assign m390 = twice_mod(m389,n); assign r390 = mult_non_zero(r389, e[389],m390) % n;
  assign m391 = twice_mod(m390,n); assign r391 = mult_non_zero(r390, e[390],m391) % n;
  assign m392 = twice_mod(m391,n); assign r392 = mult_non_zero(r391, e[391],m392) % n;
  assign m393 = twice_mod(m392,n); assign r393 = mult_non_zero(r392, e[392],m393) % n;
  assign m394 = twice_mod(m393,n); assign r394 = mult_non_zero(r393, e[393],m394) % n;
  assign m395 = twice_mod(m394,n); assign r395 = mult_non_zero(r394, e[394],m395) % n;
  assign m396 = twice_mod(m395,n); assign r396 = mult_non_zero(r395, e[395],m396) % n;
  assign m397 = twice_mod(m396,n); assign r397 = mult_non_zero(r396, e[396],m397) % n;
  assign m398 = twice_mod(m397,n); assign r398 = mult_non_zero(r397, e[397],m398) % n;
  assign m399 = twice_mod(m398,n); assign r399 = mult_non_zero(r398, e[398],m399) % n;
  assign m400 = twice_mod(m399,n); assign r400 = mult_non_zero(r399, e[399],m400) % n;
  assign m401 = twice_mod(m400,n); assign r401 = mult_non_zero(r400, e[400],m401) % n;
  assign m402 = twice_mod(m401,n); assign r402 = mult_non_zero(r401, e[401],m402) % n;
  assign m403 = twice_mod(m402,n); assign r403 = mult_non_zero(r402, e[402],m403) % n;
  assign m404 = twice_mod(m403,n); assign r404 = mult_non_zero(r403, e[403],m404) % n;
  assign m405 = twice_mod(m404,n); assign r405 = mult_non_zero(r404, e[404],m405) % n;
  assign m406 = twice_mod(m405,n); assign r406 = mult_non_zero(r405, e[405],m406) % n;
  assign m407 = twice_mod(m406,n); assign r407 = mult_non_zero(r406, e[406],m407) % n;
  assign m408 = twice_mod(m407,n); assign r408 = mult_non_zero(r407, e[407],m408) % n;
  assign m409 = twice_mod(m408,n); assign r409 = mult_non_zero(r408, e[408],m409) % n;
  assign m410 = twice_mod(m409,n); assign r410 = mult_non_zero(r409, e[409],m410) % n;
  assign m411 = twice_mod(m410,n); assign r411 = mult_non_zero(r410, e[410],m411) % n;
  assign m412 = twice_mod(m411,n); assign r412 = mult_non_zero(r411, e[411],m412) % n;
  assign m413 = twice_mod(m412,n); assign r413 = mult_non_zero(r412, e[412],m413) % n;
  assign m414 = twice_mod(m413,n); assign r414 = mult_non_zero(r413, e[413],m414) % n;
  assign m415 = twice_mod(m414,n); assign r415 = mult_non_zero(r414, e[414],m415) % n;
  assign m416 = twice_mod(m415,n); assign r416 = mult_non_zero(r415, e[415],m416) % n;
  assign m417 = twice_mod(m416,n); assign r417 = mult_non_zero(r416, e[416],m417) % n;
  assign m418 = twice_mod(m417,n); assign r418 = mult_non_zero(r417, e[417],m418) % n;
  assign m419 = twice_mod(m418,n); assign r419 = mult_non_zero(r418, e[418],m419) % n;
  assign m420 = twice_mod(m419,n); assign r420 = mult_non_zero(r419, e[419],m420) % n;
  assign m421 = twice_mod(m420,n); assign r421 = mult_non_zero(r420, e[420],m421) % n;
  assign m422 = twice_mod(m421,n); assign r422 = mult_non_zero(r421, e[421],m422) % n;
  assign m423 = twice_mod(m422,n); assign r423 = mult_non_zero(r422, e[422],m423) % n;
  assign m424 = twice_mod(m423,n); assign r424 = mult_non_zero(r423, e[423],m424) % n;
  assign m425 = twice_mod(m424,n); assign r425 = mult_non_zero(r424, e[424],m425) % n;
  assign m426 = twice_mod(m425,n); assign r426 = mult_non_zero(r425, e[425],m426) % n;
  assign m427 = twice_mod(m426,n); assign r427 = mult_non_zero(r426, e[426],m427) % n;
  assign m428 = twice_mod(m427,n); assign r428 = mult_non_zero(r427, e[427],m428) % n;
  assign m429 = twice_mod(m428,n); assign r429 = mult_non_zero(r428, e[428],m429) % n;
  assign m430 = twice_mod(m429,n); assign r430 = mult_non_zero(r429, e[429],m430) % n;
  assign m431 = twice_mod(m430,n); assign r431 = mult_non_zero(r430, e[430],m431) % n;
  assign m432 = twice_mod(m431,n); assign r432 = mult_non_zero(r431, e[431],m432) % n;
  assign m433 = twice_mod(m432,n); assign r433 = mult_non_zero(r432, e[432],m433) % n;
  assign m434 = twice_mod(m433,n); assign r434 = mult_non_zero(r433, e[433],m434) % n;
  assign m435 = twice_mod(m434,n); assign r435 = mult_non_zero(r434, e[434],m435) % n;
  assign m436 = twice_mod(m435,n); assign r436 = mult_non_zero(r435, e[435],m436) % n;
  assign m437 = twice_mod(m436,n); assign r437 = mult_non_zero(r436, e[436],m437) % n;
  assign m438 = twice_mod(m437,n); assign r438 = mult_non_zero(r437, e[437],m438) % n;
  assign m439 = twice_mod(m438,n); assign r439 = mult_non_zero(r438, e[438],m439) % n;
  assign m440 = twice_mod(m439,n); assign r440 = mult_non_zero(r439, e[439],m440) % n;
  assign m441 = twice_mod(m440,n); assign r441 = mult_non_zero(r440, e[440],m441) % n;
  assign m442 = twice_mod(m441,n); assign r442 = mult_non_zero(r441, e[441],m442) % n;
  assign m443 = twice_mod(m442,n); assign r443 = mult_non_zero(r442, e[442],m443) % n;
  assign m444 = twice_mod(m443,n); assign r444 = mult_non_zero(r443, e[443],m444) % n;
  assign m445 = twice_mod(m444,n); assign r445 = mult_non_zero(r444, e[444],m445) % n;
  assign m446 = twice_mod(m445,n); assign r446 = mult_non_zero(r445, e[445],m446) % n;
  assign m447 = twice_mod(m446,n); assign r447 = mult_non_zero(r446, e[446],m447) % n;
  assign m448 = twice_mod(m447,n); assign r448 = mult_non_zero(r447, e[447],m448) % n;
  assign m449 = twice_mod(m448,n); assign r449 = mult_non_zero(r448, e[448],m449) % n;
  assign m450 = twice_mod(m449,n); assign r450 = mult_non_zero(r449, e[449],m450) % n;
  assign m451 = twice_mod(m450,n); assign r451 = mult_non_zero(r450, e[450],m451) % n;
  assign m452 = twice_mod(m451,n); assign r452 = mult_non_zero(r451, e[451],m452) % n;
  assign m453 = twice_mod(m452,n); assign r453 = mult_non_zero(r452, e[452],m453) % n;
  assign m454 = twice_mod(m453,n); assign r454 = mult_non_zero(r453, e[453],m454) % n;
  assign m455 = twice_mod(m454,n); assign r455 = mult_non_zero(r454, e[454],m455) % n;
  assign m456 = twice_mod(m455,n); assign r456 = mult_non_zero(r455, e[455],m456) % n;
  assign m457 = twice_mod(m456,n); assign r457 = mult_non_zero(r456, e[456],m457) % n;
  assign m458 = twice_mod(m457,n); assign r458 = mult_non_zero(r457, e[457],m458) % n;
  assign m459 = twice_mod(m458,n); assign r459 = mult_non_zero(r458, e[458],m459) % n;
  assign m460 = twice_mod(m459,n); assign r460 = mult_non_zero(r459, e[459],m460) % n;
  assign m461 = twice_mod(m460,n); assign r461 = mult_non_zero(r460, e[460],m461) % n;
  assign m462 = twice_mod(m461,n); assign r462 = mult_non_zero(r461, e[461],m462) % n;
  assign m463 = twice_mod(m462,n); assign r463 = mult_non_zero(r462, e[462],m463) % n;
  assign m464 = twice_mod(m463,n); assign r464 = mult_non_zero(r463, e[463],m464) % n;
  assign m465 = twice_mod(m464,n); assign r465 = mult_non_zero(r464, e[464],m465) % n;
  assign m466 = twice_mod(m465,n); assign r466 = mult_non_zero(r465, e[465],m466) % n;
  assign m467 = twice_mod(m466,n); assign r467 = mult_non_zero(r466, e[466],m467) % n;
  assign m468 = twice_mod(m467,n); assign r468 = mult_non_zero(r467, e[467],m468) % n;
  assign m469 = twice_mod(m468,n); assign r469 = mult_non_zero(r468, e[468],m469) % n;
  assign m470 = twice_mod(m469,n); assign r470 = mult_non_zero(r469, e[469],m470) % n;
  assign m471 = twice_mod(m470,n); assign r471 = mult_non_zero(r470, e[470],m471) % n;
  assign m472 = twice_mod(m471,n); assign r472 = mult_non_zero(r471, e[471],m472) % n;
  assign m473 = twice_mod(m472,n); assign r473 = mult_non_zero(r472, e[472],m473) % n;
  assign m474 = twice_mod(m473,n); assign r474 = mult_non_zero(r473, e[473],m474) % n;
  assign m475 = twice_mod(m474,n); assign r475 = mult_non_zero(r474, e[474],m475) % n;
  assign m476 = twice_mod(m475,n); assign r476 = mult_non_zero(r475, e[475],m476) % n;
  assign m477 = twice_mod(m476,n); assign r477 = mult_non_zero(r476, e[476],m477) % n;
  assign m478 = twice_mod(m477,n); assign r478 = mult_non_zero(r477, e[477],m478) % n;
  assign m479 = twice_mod(m478,n); assign r479 = mult_non_zero(r478, e[478],m479) % n;
  assign m480 = twice_mod(m479,n); assign r480 = mult_non_zero(r479, e[479],m480) % n;
  assign m481 = twice_mod(m480,n); assign r481 = mult_non_zero(r480, e[480],m481) % n;
  assign m482 = twice_mod(m481,n); assign r482 = mult_non_zero(r481, e[481],m482) % n;
  assign m483 = twice_mod(m482,n); assign r483 = mult_non_zero(r482, e[482],m483) % n;
  assign m484 = twice_mod(m483,n); assign r484 = mult_non_zero(r483, e[483],m484) % n;
  assign m485 = twice_mod(m484,n); assign r485 = mult_non_zero(r484, e[484],m485) % n;
  assign m486 = twice_mod(m485,n); assign r486 = mult_non_zero(r485, e[485],m486) % n;
  assign m487 = twice_mod(m486,n); assign r487 = mult_non_zero(r486, e[486],m487) % n;
  assign m488 = twice_mod(m487,n); assign r488 = mult_non_zero(r487, e[487],m488) % n;
  assign m489 = twice_mod(m488,n); assign r489 = mult_non_zero(r488, e[488],m489) % n;
  assign m490 = twice_mod(m489,n); assign r490 = mult_non_zero(r489, e[489],m490) % n;
  assign m491 = twice_mod(m490,n); assign r491 = mult_non_zero(r490, e[490],m491) % n;
  assign m492 = twice_mod(m491,n); assign r492 = mult_non_zero(r491, e[491],m492) % n;
  assign m493 = twice_mod(m492,n); assign r493 = mult_non_zero(r492, e[492],m493) % n;
  assign m494 = twice_mod(m493,n); assign r494 = mult_non_zero(r493, e[493],m494) % n;
  assign m495 = twice_mod(m494,n); assign r495 = mult_non_zero(r494, e[494],m495) % n;
  assign m496 = twice_mod(m495,n); assign r496 = mult_non_zero(r495, e[495],m496) % n;
  assign m497 = twice_mod(m496,n); assign r497 = mult_non_zero(r496, e[496],m497) % n;
  assign m498 = twice_mod(m497,n); assign r498 = mult_non_zero(r497, e[497],m498) % n;
  assign m499 = twice_mod(m498,n); assign r499 = mult_non_zero(r498, e[498],m499) % n;
  assign m500 = twice_mod(m499,n); assign r500 = mult_non_zero(r499, e[499],m500) % n;
  assign m501 = twice_mod(m500,n); assign r501 = mult_non_zero(r500, e[500],m501) % n;
  assign m502 = twice_mod(m501,n); assign r502 = mult_non_zero(r501, e[501],m502) % n;
  assign m503 = twice_mod(m502,n); assign r503 = mult_non_zero(r502, e[502],m503) % n;
  assign m504 = twice_mod(m503,n); assign r504 = mult_non_zero(r503, e[503],m504) % n;
  assign m505 = twice_mod(m504,n); assign r505 = mult_non_zero(r504, e[504],m505) % n;
  assign m506 = twice_mod(m505,n); assign r506 = mult_non_zero(r505, e[505],m506) % n;
  assign m507 = twice_mod(m506,n); assign r507 = mult_non_zero(r506, e[506],m507) % n;
  assign m508 = twice_mod(m507,n); assign r508 = mult_non_zero(r507, e[507],m508) % n;
  assign m509 = twice_mod(m508,n); assign r509 = mult_non_zero(r508, e[508],m509) % n;
  assign m510 = twice_mod(m509,n); assign r510 = mult_non_zero(r509, e[509],m510) % n;
  assign m511 = twice_mod(m510,n); assign r511 = mult_non_zero(r510, e[510],m511) % n;
  assign m512 = twice_mod(m511,n); assign r512 = mult_non_zero(r511, e[511],m512) % n;

  assign r = r512;

  function [1023:0] mult;
    input [511:0] m,n;
    mult = m * n;
  endfunction

  function [1023:0] mult_non_zero;
    input [511:0] r;
    input [1:0]   b;
    input [511:0] m;
    mult_non_zero = mult(r , (b == 1'b1 ? m : 1) );
  endfunction

  function [511:0] twice_mod;
    input [511:0] m, n;
    twice_mod = mult(m,m) % n;
  endfunction

endmodule





module test;
  reg  [0:511]e,n,m;
  wire [0:511]r;

  initial begin
      n  <= 16;
      m  <= 3;
      e  <= 3;
    #1
      n  <= 1024;
      m  <= 8;
      e  <= 2;
    #1
      n  <= 512'hA940A3603B2A227D3B7E945F528E92214A4F3DDAED3411A669E34AF64D59302BFAF333F281AF17C483901AF2490BC8AD3827ED7AC03A97A7B446C6AF84D2803B;
      m  <= 512'h166cc193544bf5666277170104384363562a8ff3c25ffb93f7c49244eb55ad654f51da4bbca25fa5f3fe727dbecdd0659af3d1b7b6ac8035d6cab2576aee4ce8;
      e  <= 512'h10001;
      // r:3030303030303030303030303030303030303030303030303030303030303030303030303030303030303030303030303030303030303030303030303030300a
  end

  modexp1 modexp(e,n,m,r);

  initial begin
    $monitor ($stime , " hello world e:%h n:%h m:%h r:%h ",e,n,m,r);
//    $monitor ($stime , " r001 %h r002 %h r003 %h",modexp.r001,modexp.r002,modexp.r003);
//    $monitor ($stime , " m001 %h m002 %h m003 %h",modexp.m001,modexp.m002,modexp.m003);
//    $monitor ($stime , " e[1] %h e[2] %h e[3] %h",modexp.e[0],modexp.e[1],modexp.e[2]);
  end

endmodule
