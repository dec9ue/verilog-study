

module modexp1 ( e ,n,m, r);
  input[511:0] e,n,m;
  output[511:0] r;

  wire [511:0] m000, r000; wire [511:0] m001, r001; wire [511:0] m002, r002; wire [511:0] m003, r003; wire [511:0] m004, r004; wire [511:0] m005, r005; wire [511:0] m006, r006; wire [511:0] m007, r007; wire [511:0] m008, r008; wire [511:0] m009, r009; wire [511:0] m010, r010; wire [511:0] m011, r011; wire [511:0] m012, r012; wire [511:0] m013, r013; wire [511:0] m014, r014; wire [511:0] m015, r015; wire [511:0] m016, r016; wire [511:0] m017, r017; wire [511:0] m018, r018; wire [511:0] m019, r019; wire [511:0] m020, r020; wire [511:0] m021, r021; wire [511:0] m022, r022; wire [511:0] m023, r023; wire [511:0] m024, r024; wire [511:0] m025, r025; wire [511:0] m026, r026; wire [511:0] m027, r027; wire [511:0] m028, r028; wire [511:0] m029, r029; wire [511:0] m030, r030; wire [511:0] m031, r031; wire [511:0] m032, r032; wire [511:0] m033, r033; wire [511:0] m034, r034; wire [511:0] m035, r035; wire [511:0] m036, r036; wire [511:0] m037, r037; wire [511:0] m038, r038; wire [511:0] m039, r039; wire [511:0] m040, r040; wire [511:0] m041, r041; wire [511:0] m042, r042; wire [511:0] m043, r043; wire [511:0] m044, r044; wire [511:0] m045, r045; wire [511:0] m046, r046; wire [511:0] m047, r047; wire [511:0] m048, r048; wire [511:0] m049, r049; wire [511:0] m050, r050; wire [511:0] m051, r051; wire [511:0] m052, r052; wire [511:0] m053, r053; wire [511:0] m054, r054; wire [511:0] m055, r055; wire [511:0] m056, r056; wire [511:0] m057, r057; wire [511:0] m058, r058; wire [511:0] m059, r059; wire [511:0] m060, r060; wire [511:0] m061, r061; wire [511:0] m062, r062; wire [511:0] m063, r063; wire [511:0] m064, r064; wire [511:0] m065, r065; wire [511:0] m066, r066; wire [511:0] m067, r067; wire [511:0] m068, r068; wire [511:0] m069, r069; wire [511:0] m070, r070; wire [511:0] m071, r071; wire [511:0] m072, r072; wire [511:0] m073, r073; wire [511:0] m074, r074; wire [511:0] m075, r075; wire [511:0] m076, r076; wire [511:0] m077, r077; wire [511:0] m078, r078; wire [511:0] m079, r079; wire [511:0] m080, r080; wire [511:0] m081, r081; wire [511:0] m082, r082; wire [511:0] m083, r083; wire [511:0] m084, r084; wire [511:0] m085, r085; wire [511:0] m086, r086; wire [511:0] m087, r087; wire [511:0] m088, r088; wire [511:0] m089, r089; wire [511:0] m090, r090; wire [511:0] m091, r091; wire [511:0] m092, r092; wire [511:0] m093, r093; wire [511:0] m094, r094; wire [511:0] m095, r095; wire [511:0] m096, r096; wire [511:0] m097, r097; wire [511:0] m098, r098; wire [511:0] m099, r099; wire [511:0] m100, r100; wire [511:0] m101, r101; wire [511:0] m102, r102; wire [511:0] m103, r103; wire [511:0] m104, r104; wire [511:0] m105, r105; wire [511:0] m106, r106; wire [511:0] m107, r107; wire [511:0] m108, r108; wire [511:0] m109, r109; wire [511:0] m110, r110; wire [511:0] m111, r111; wire [511:0] m112, r112; wire [511:0] m113, r113; wire [511:0] m114, r114; wire [511:0] m115, r115; wire [511:0] m116, r116; wire [511:0] m117, r117; wire [511:0] m118, r118; wire [511:0] m119, r119; wire [511:0] m120, r120; wire [511:0] m121, r121; wire [511:0] m122, r122; wire [511:0] m123, r123; wire [511:0] m124, r124; wire [511:0] m125, r125; wire [511:0] m126, r126; wire [511:0] m127, r127;
  wire [511:0] m128, r128; wire [511:0] m129, r129; wire [511:0] m130, r130; wire [511:0] m131, r131; wire [511:0] m132, r132; wire [511:0] m133, r133; wire [511:0] m134, r134; wire [511:0] m135, r135; wire [511:0] m136, r136; wire [511:0] m137, r137; wire [511:0] m138, r138; wire [511:0] m139, r139; wire [511:0] m140, r140; wire [511:0] m141, r141; wire [511:0] m142, r142; wire [511:0] m143, r143; wire [511:0] m144, r144; wire [511:0] m145, r145; wire [511:0] m146, r146; wire [511:0] m147, r147; wire [511:0] m148, r148; wire [511:0] m149, r149; wire [511:0] m150, r150; wire [511:0] m151, r151; wire [511:0] m152, r152; wire [511:0] m153, r153; wire [511:0] m154, r154; wire [511:0] m155, r155; wire [511:0] m156, r156; wire [511:0] m157, r157; wire [511:0] m158, r158; wire [511:0] m159, r159; wire [511:0] m160, r160; wire [511:0] m161, r161; wire [511:0] m162, r162; wire [511:0] m163, r163; wire [511:0] m164, r164; wire [511:0] m165, r165; wire [511:0] m166, r166; wire [511:0] m167, r167; wire [511:0] m168, r168; wire [511:0] m169, r169; wire [511:0] m170, r170; wire [511:0] m171, r171; wire [511:0] m172, r172; wire [511:0] m173, r173; wire [511:0] m174, r174; wire [511:0] m175, r175; wire [511:0] m176, r176; wire [511:0] m177, r177; wire [511:0] m178, r178; wire [511:0] m179, r179; wire [511:0] m180, r180; wire [511:0] m181, r181; wire [511:0] m182, r182; wire [511:0] m183, r183; wire [511:0] m184, r184; wire [511:0] m185, r185; wire [511:0] m186, r186; wire [511:0] m187, r187; wire [511:0] m188, r188; wire [511:0] m189, r189; wire [511:0] m190, r190; wire [511:0] m191, r191; wire [511:0] m192, r192; wire [511:0] m193, r193; wire [511:0] m194, r194; wire [511:0] m195, r195; wire [511:0] m196, r196; wire [511:0] m197, r197; wire [511:0] m198, r198; wire [511:0] m199, r199; wire [511:0] m200, r200; wire [511:0] m201, r201; wire [511:0] m202, r202; wire [511:0] m203, r203; wire [511:0] m204, r204; wire [511:0] m205, r205; wire [511:0] m206, r206; wire [511:0] m207, r207; wire [511:0] m208, r208; wire [511:0] m209, r209; wire [511:0] m210, r210; wire [511:0] m211, r211; wire [511:0] m212, r212; wire [511:0] m213, r213; wire [511:0] m214, r214; wire [511:0] m215, r215; wire [511:0] m216, r216; wire [511:0] m217, r217; wire [511:0] m218, r218; wire [511:0] m219, r219; wire [511:0] m220, r220; wire [511:0] m221, r221; wire [511:0] m222, r222; wire [511:0] m223, r223; wire [511:0] m224, r224; wire [511:0] m225, r225; wire [511:0] m226, r226; wire [511:0] m227, r227; wire [511:0] m228, r228; wire [511:0] m229, r229; wire [511:0] m230, r230; wire [511:0] m231, r231; wire [511:0] m232, r232; wire [511:0] m233, r233; wire [511:0] m234, r234; wire [511:0] m235, r235; wire [511:0] m236, r236; wire [511:0] m237, r237; wire [511:0] m238, r238; wire [511:0] m239, r239; wire [511:0] m240, r240; wire [511:0] m241, r241; wire [511:0] m242, r242; wire [511:0] m243, r243; wire [511:0] m244, r244; wire [511:0] m245, r245; wire [511:0] m246, r246; wire [511:0] m247, r247; wire [511:0] m248, r248; wire [511:0] m249, r249; wire [511:0] m250, r250; wire [511:0] m251, r251; wire [511:0] m252, r252; wire [511:0] m253, r253; wire [511:0] m254, r254; wire [511:0] m255, r255;
  wire [511:0] m256, r256; wire [511:0] m257, r257; wire [511:0] m258, r258; wire [511:0] m259, r259; wire [511:0] m260, r260; wire [511:0] m261, r261; wire [511:0] m262, r262; wire [511:0] m263, r263; wire [511:0] m264, r264; wire [511:0] m265, r265; wire [511:0] m266, r266; wire [511:0] m267, r267; wire [511:0] m268, r268; wire [511:0] m269, r269; wire [511:0] m270, r270; wire [511:0] m271, r271; wire [511:0] m272, r272; wire [511:0] m273, r273; wire [511:0] m274, r274; wire [511:0] m275, r275; wire [511:0] m276, r276; wire [511:0] m277, r277; wire [511:0] m278, r278; wire [511:0] m279, r279; wire [511:0] m280, r280; wire [511:0] m281, r281; wire [511:0] m282, r282; wire [511:0] m283, r283; wire [511:0] m284, r284; wire [511:0] m285, r285; wire [511:0] m286, r286; wire [511:0] m287, r287; wire [511:0] m288, r288; wire [511:0] m289, r289; wire [511:0] m290, r290; wire [511:0] m291, r291; wire [511:0] m292, r292; wire [511:0] m293, r293; wire [511:0] m294, r294; wire [511:0] m295, r295; wire [511:0] m296, r296; wire [511:0] m297, r297; wire [511:0] m298, r298; wire [511:0] m299, r299; wire [511:0] m300, r300; wire [511:0] m301, r301; wire [511:0] m302, r302; wire [511:0] m303, r303; wire [511:0] m304, r304; wire [511:0] m305, r305; wire [511:0] m306, r306; wire [511:0] m307, r307; wire [511:0] m308, r308; wire [511:0] m309, r309; wire [511:0] m310, r310; wire [511:0] m311, r311; wire [511:0] m312, r312; wire [511:0] m313, r313; wire [511:0] m314, r314; wire [511:0] m315, r315; wire [511:0] m316, r316; wire [511:0] m317, r317; wire [511:0] m318, r318; wire [511:0] m319, r319; wire [511:0] m320, r320; wire [511:0] m321, r321; wire [511:0] m322, r322; wire [511:0] m323, r323; wire [511:0] m324, r324; wire [511:0] m325, r325; wire [511:0] m326, r326; wire [511:0] m327, r327; wire [511:0] m328, r328; wire [511:0] m329, r329; wire [511:0] m330, r330; wire [511:0] m331, r331; wire [511:0] m332, r332; wire [511:0] m333, r333; wire [511:0] m334, r334; wire [511:0] m335, r335; wire [511:0] m336, r336; wire [511:0] m337, r337; wire [511:0] m338, r338; wire [511:0] m339, r339; wire [511:0] m340, r340; wire [511:0] m341, r341; wire [511:0] m342, r342; wire [511:0] m343, r343; wire [511:0] m344, r344; wire [511:0] m345, r345; wire [511:0] m346, r346; wire [511:0] m347, r347; wire [511:0] m348, r348; wire [511:0] m349, r349; wire [511:0] m350, r350; wire [511:0] m351, r351; wire [511:0] m352, r352; wire [511:0] m353, r353; wire [511:0] m354, r354; wire [511:0] m355, r355; wire [511:0] m356, r356; wire [511:0] m357, r357; wire [511:0] m358, r358; wire [511:0] m359, r359; wire [511:0] m360, r360; wire [511:0] m361, r361; wire [511:0] m362, r362; wire [511:0] m363, r363; wire [511:0] m364, r364; wire [511:0] m365, r365; wire [511:0] m366, r366; wire [511:0] m367, r367; wire [511:0] m368, r368; wire [511:0] m369, r369; wire [511:0] m370, r370; wire [511:0] m371, r371; wire [511:0] m372, r372; wire [511:0] m373, r373; wire [511:0] m374, r374; wire [511:0] m375, r375; wire [511:0] m376, r376; wire [511:0] m377, r377; wire [511:0] m378, r378; wire [511:0] m379, r379; wire [511:0] m380, r380; wire [511:0] m381, r381; wire [511:0] m382, r382; wire [511:0] m383, r383;
  wire [511:0] m384, r384; wire [511:0] m385, r385; wire [511:0] m386, r386; wire [511:0] m387, r387; wire [511:0] m388, r388; wire [511:0] m389, r389; wire [511:0] m390, r390; wire [511:0] m391, r391; wire [511:0] m392, r392; wire [511:0] m393, r393; wire [511:0] m394, r394; wire [511:0] m395, r395; wire [511:0] m396, r396; wire [511:0] m397, r397; wire [511:0] m398, r398; wire [511:0] m399, r399; wire [511:0] m400, r400; wire [511:0] m401, r401; wire [511:0] m402, r402; wire [511:0] m403, r403; wire [511:0] m404, r404; wire [511:0] m405, r405; wire [511:0] m406, r406; wire [511:0] m407, r407; wire [511:0] m408, r408; wire [511:0] m409, r409; wire [511:0] m410, r410; wire [511:0] m411, r411; wire [511:0] m412, r412; wire [511:0] m413, r413; wire [511:0] m414, r414; wire [511:0] m415, r415; wire [511:0] m416, r416; wire [511:0] m417, r417; wire [511:0] m418, r418; wire [511:0] m419, r419; wire [511:0] m420, r420; wire [511:0] m421, r421; wire [511:0] m422, r422; wire [511:0] m423, r423; wire [511:0] m424, r424; wire [511:0] m425, r425; wire [511:0] m426, r426; wire [511:0] m427, r427; wire [511:0] m428, r428; wire [511:0] m429, r429; wire [511:0] m430, r430; wire [511:0] m431, r431; wire [511:0] m432, r432; wire [511:0] m433, r433; wire [511:0] m434, r434; wire [511:0] m435, r435; wire [511:0] m436, r436; wire [511:0] m437, r437; wire [511:0] m438, r438; wire [511:0] m439, r439; wire [511:0] m440, r440; wire [511:0] m441, r441; wire [511:0] m442, r442; wire [511:0] m443, r443; wire [511:0] m444, r444; wire [511:0] m445, r445; wire [511:0] m446, r446; wire [511:0] m447, r447; wire [511:0] m448, r448; wire [511:0] m449, r449; wire [511:0] m450, r450; wire [511:0] m451, r451; wire [511:0] m452, r452; wire [511:0] m453, r453; wire [511:0] m454, r454; wire [511:0] m455, r455; wire [511:0] m456, r456; wire [511:0] m457, r457; wire [511:0] m458, r458; wire [511:0] m459, r459; wire [511:0] m460, r460; wire [511:0] m461, r461; wire [511:0] m462, r462; wire [511:0] m463, r463; wire [511:0] m464, r464; wire [511:0] m465, r465; wire [511:0] m466, r466; wire [511:0] m467, r467; wire [511:0] m468, r468; wire [511:0] m469, r469; wire [511:0] m470, r470; wire [511:0] m471, r471; wire [511:0] m472, r472; wire [511:0] m473, r473; wire [511:0] m474, r474; wire [511:0] m475, r475; wire [511:0] m476, r476; wire [511:0] m477, r477; wire [511:0] m478, r478; wire [511:0] m479, r479; wire [511:0] m480, r480; wire [511:0] m481, r481; wire [511:0] m482, r482; wire [511:0] m483, r483; wire [511:0] m484, r484; wire [511:0] m485, r485; wire [511:0] m486, r486; wire [511:0] m487, r487; wire [511:0] m488, r488; wire [511:0] m489, r489; wire [511:0] m490, r490; wire [511:0] m491, r491; wire [511:0] m492, r492; wire [511:0] m493, r493; wire [511:0] m494, r494; wire [511:0] m495, r495; wire [511:0] m496, r496; wire [511:0] m497, r497; wire [511:0] m498, r498; wire [511:0] m499, r499; wire [511:0] m500, r500; wire [511:0] m501, r501; wire [511:0] m502, r502; wire [511:0] m503, r503; wire [511:0] m504, r504; wire [511:0] m505, r505; wire [511:0] m506, r506; wire [511:0] m507, r507; wire [511:0] m508, r508; wire [511:0] m509, r509; wire [511:0] m510, r510; wire [511:0] m511, r511;
  wire [511:0] m512, r512;

  assign m001 = m;
  assign r001 = (1 * (1 + e[0] * (m001 - 1))) % n;

  assign m002 = twice_mod(m001,n); assign r002 = (r001 * (1+ e[1] * (m002 - 1))) % n;
  assign m003 = twice_mod(m002,n); assign r003 = (r002 * (1+ e[2] * (m003 - 1))) % n;
  assign m004 = twice_mod(m003,n); assign r004 = (r003 * (1+ e[3] * (m004 - 1))) % n;
  assign m005 = twice_mod(m004,n); assign r005 = (r004 * (1+ e[4] * (m005 - 1))) % n;
  assign m006 = twice_mod(m005,n); assign r006 = (r005 * (1+ e[5] * (m006 - 1))) % n;
  assign m007 = twice_mod(m006,n); assign r007 = (r006 * (1+ e[6] * (m007 - 1))) % n;
  assign m008 = twice_mod(m007,n); assign r008 = (r007 * (1+ e[7] * (m008 - 1))) % n;
  assign m009 = twice_mod(m008,n); assign r009 = (r008 * (1+ e[8] * (m009 - 1))) % n;
  assign m010 = twice_mod(m009,n); assign r010 = (r009 * (1+ e[9] * (m010 - 1))) % n;
  assign m011 = twice_mod(m010,n); assign r011 = (r010 * (1+ e[10] * (m011 - 1))) % n;
  assign m012 = twice_mod(m011,n); assign r012 = (r011 * (1+ e[11] * (m012 - 1))) % n;
  assign m013 = twice_mod(m012,n); assign r013 = (r012 * (1+ e[12] * (m013 - 1))) % n;
  assign m014 = twice_mod(m013,n); assign r014 = (r013 * (1+ e[13] * (m014 - 1))) % n;
  assign m015 = twice_mod(m014,n); assign r015 = (r014 * (1+ e[14] * (m015 - 1))) % n;
  assign m016 = twice_mod(m015,n); assign r016 = (r015 * (1+ e[15] * (m016 - 1))) % n;
  assign m017 = twice_mod(m016,n); assign r017 = (r016 * (1+ e[16] * (m017 - 1))) % n;
  assign m018 = twice_mod(m017,n); assign r018 = (r017 * (1+ e[17] * (m018 - 1))) % n;
  assign m019 = twice_mod(m018,n); assign r019 = (r018 * (1+ e[18] * (m019 - 1))) % n;
  assign m020 = twice_mod(m019,n); assign r020 = (r019 * (1+ e[19] * (m020 - 1))) % n;
  assign m021 = twice_mod(m020,n); assign r021 = (r020 * (1+ e[20] * (m021 - 1))) % n;
  assign m022 = twice_mod(m021,n); assign r022 = (r021 * (1+ e[21] * (m022 - 1))) % n;
  assign m023 = twice_mod(m022,n); assign r023 = (r022 * (1+ e[22] * (m023 - 1))) % n;
  assign m024 = twice_mod(m023,n); assign r024 = (r023 * (1+ e[23] * (m024 - 1))) % n;
  assign m025 = twice_mod(m024,n); assign r025 = (r024 * (1+ e[24] * (m025 - 1))) % n;
  assign m026 = twice_mod(m025,n); assign r026 = (r025 * (1+ e[25] * (m026 - 1))) % n;
  assign m027 = twice_mod(m026,n); assign r027 = (r026 * (1+ e[26] * (m027 - 1))) % n;
  assign m028 = twice_mod(m027,n); assign r028 = (r027 * (1+ e[27] * (m028 - 1))) % n;
  assign m029 = twice_mod(m028,n); assign r029 = (r028 * (1+ e[28] * (m029 - 1))) % n;
  assign m030 = twice_mod(m029,n); assign r030 = (r029 * (1+ e[29] * (m030 - 1))) % n;
  assign m031 = twice_mod(m030,n); assign r031 = (r030 * (1+ e[30] * (m031 - 1))) % n;
  assign m032 = twice_mod(m031,n); assign r032 = (r031 * (1+ e[31] * (m032 - 1))) % n;
  assign m033 = twice_mod(m032,n); assign r033 = (r032 * (1+ e[32] * (m033 - 1))) % n;
  assign m034 = twice_mod(m033,n); assign r034 = (r033 * (1+ e[33] * (m034 - 1))) % n;
  assign m035 = twice_mod(m034,n); assign r035 = (r034 * (1+ e[34] * (m035 - 1))) % n;
  assign m036 = twice_mod(m035,n); assign r036 = (r035 * (1+ e[35] * (m036 - 1))) % n;
  assign m037 = twice_mod(m036,n); assign r037 = (r036 * (1+ e[36] * (m037 - 1))) % n;
  assign m038 = twice_mod(m037,n); assign r038 = (r037 * (1+ e[37] * (m038 - 1))) % n;
  assign m039 = twice_mod(m038,n); assign r039 = (r038 * (1+ e[38] * (m039 - 1))) % n;
  assign m040 = twice_mod(m039,n); assign r040 = (r039 * (1+ e[39] * (m040 - 1))) % n;
  assign m041 = twice_mod(m040,n); assign r041 = (r040 * (1+ e[40] * (m041 - 1))) % n;
  assign m042 = twice_mod(m041,n); assign r042 = (r041 * (1+ e[41] * (m042 - 1))) % n;
  assign m043 = twice_mod(m042,n); assign r043 = (r042 * (1+ e[42] * (m043 - 1))) % n;
  assign m044 = twice_mod(m043,n); assign r044 = (r043 * (1+ e[43] * (m044 - 1))) % n;
  assign m045 = twice_mod(m044,n); assign r045 = (r044 * (1+ e[44] * (m045 - 1))) % n;
  assign m046 = twice_mod(m045,n); assign r046 = (r045 * (1+ e[45] * (m046 - 1))) % n;
  assign m047 = twice_mod(m046,n); assign r047 = (r046 * (1+ e[46] * (m047 - 1))) % n;
  assign m048 = twice_mod(m047,n); assign r048 = (r047 * (1+ e[47] * (m048 - 1))) % n;
  assign m049 = twice_mod(m048,n); assign r049 = (r048 * (1+ e[48] * (m049 - 1))) % n;
  assign m050 = twice_mod(m049,n); assign r050 = (r049 * (1+ e[49] * (m050 - 1))) % n;
  assign m051 = twice_mod(m050,n); assign r051 = (r050 * (1+ e[50] * (m051 - 1))) % n;
  assign m052 = twice_mod(m051,n); assign r052 = (r051 * (1+ e[51] * (m052 - 1))) % n;
  assign m053 = twice_mod(m052,n); assign r053 = (r052 * (1+ e[52] * (m053 - 1))) % n;
  assign m054 = twice_mod(m053,n); assign r054 = (r053 * (1+ e[53] * (m054 - 1))) % n;
  assign m055 = twice_mod(m054,n); assign r055 = (r054 * (1+ e[54] * (m055 - 1))) % n;
  assign m056 = twice_mod(m055,n); assign r056 = (r055 * (1+ e[55] * (m056 - 1))) % n;
  assign m057 = twice_mod(m056,n); assign r057 = (r056 * (1+ e[56] * (m057 - 1))) % n;
  assign m058 = twice_mod(m057,n); assign r058 = (r057 * (1+ e[57] * (m058 - 1))) % n;
  assign m059 = twice_mod(m058,n); assign r059 = (r058 * (1+ e[58] * (m059 - 1))) % n;
  assign m060 = twice_mod(m059,n); assign r060 = (r059 * (1+ e[59] * (m060 - 1))) % n;
  assign m061 = twice_mod(m060,n); assign r061 = (r060 * (1+ e[60] * (m061 - 1))) % n;
  assign m062 = twice_mod(m061,n); assign r062 = (r061 * (1+ e[61] * (m062 - 1))) % n;
  assign m063 = twice_mod(m062,n); assign r063 = (r062 * (1+ e[62] * (m063 - 1))) % n;
  assign m064 = twice_mod(m063,n); assign r064 = (r063 * (1+ e[63] * (m064 - 1))) % n;
  assign m065 = twice_mod(m064,n); assign r065 = (r064 * (1+ e[64] * (m065 - 1))) % n;
  assign m066 = twice_mod(m065,n); assign r066 = (r065 * (1+ e[65] * (m066 - 1))) % n;
  assign m067 = twice_mod(m066,n); assign r067 = (r066 * (1+ e[66] * (m067 - 1))) % n;
  assign m068 = twice_mod(m067,n); assign r068 = (r067 * (1+ e[67] * (m068 - 1))) % n;
  assign m069 = twice_mod(m068,n); assign r069 = (r068 * (1+ e[68] * (m069 - 1))) % n;
  assign m070 = twice_mod(m069,n); assign r070 = (r069 * (1+ e[69] * (m070 - 1))) % n;
  assign m071 = twice_mod(m070,n); assign r071 = (r070 * (1+ e[70] * (m071 - 1))) % n;
  assign m072 = twice_mod(m071,n); assign r072 = (r071 * (1+ e[71] * (m072 - 1))) % n;
  assign m073 = twice_mod(m072,n); assign r073 = (r072 * (1+ e[72] * (m073 - 1))) % n;
  assign m074 = twice_mod(m073,n); assign r074 = (r073 * (1+ e[73] * (m074 - 1))) % n;
  assign m075 = twice_mod(m074,n); assign r075 = (r074 * (1+ e[74] * (m075 - 1))) % n;
  assign m076 = twice_mod(m075,n); assign r076 = (r075 * (1+ e[75] * (m076 - 1))) % n;
  assign m077 = twice_mod(m076,n); assign r077 = (r076 * (1+ e[76] * (m077 - 1))) % n;
  assign m078 = twice_mod(m077,n); assign r078 = (r077 * (1+ e[77] * (m078 - 1))) % n;
  assign m079 = twice_mod(m078,n); assign r079 = (r078 * (1+ e[78] * (m079 - 1))) % n;
  assign m080 = twice_mod(m079,n); assign r080 = (r079 * (1+ e[79] * (m080 - 1))) % n;
  assign m081 = twice_mod(m080,n); assign r081 = (r080 * (1+ e[80] * (m081 - 1))) % n;
  assign m082 = twice_mod(m081,n); assign r082 = (r081 * (1+ e[81] * (m082 - 1))) % n;
  assign m083 = twice_mod(m082,n); assign r083 = (r082 * (1+ e[82] * (m083 - 1))) % n;
  assign m084 = twice_mod(m083,n); assign r084 = (r083 * (1+ e[83] * (m084 - 1))) % n;
  assign m085 = twice_mod(m084,n); assign r085 = (r084 * (1+ e[84] * (m085 - 1))) % n;
  assign m086 = twice_mod(m085,n); assign r086 = (r085 * (1+ e[85] * (m086 - 1))) % n;
  assign m087 = twice_mod(m086,n); assign r087 = (r086 * (1+ e[86] * (m087 - 1))) % n;
  assign m088 = twice_mod(m087,n); assign r088 = (r087 * (1+ e[87] * (m088 - 1))) % n;
  assign m089 = twice_mod(m088,n); assign r089 = (r088 * (1+ e[88] * (m089 - 1))) % n;
  assign m090 = twice_mod(m089,n); assign r090 = (r089 * (1+ e[89] * (m090 - 1))) % n;
  assign m091 = twice_mod(m090,n); assign r091 = (r090 * (1+ e[90] * (m091 - 1))) % n;
  assign m092 = twice_mod(m091,n); assign r092 = (r091 * (1+ e[91] * (m092 - 1))) % n;
  assign m093 = twice_mod(m092,n); assign r093 = (r092 * (1+ e[92] * (m093 - 1))) % n;
  assign m094 = twice_mod(m093,n); assign r094 = (r093 * (1+ e[93] * (m094 - 1))) % n;
  assign m095 = twice_mod(m094,n); assign r095 = (r094 * (1+ e[94] * (m095 - 1))) % n;
  assign m096 = twice_mod(m095,n); assign r096 = (r095 * (1+ e[95] * (m096 - 1))) % n;
  assign m097 = twice_mod(m096,n); assign r097 = (r096 * (1+ e[96] * (m097 - 1))) % n;
  assign m098 = twice_mod(m097,n); assign r098 = (r097 * (1+ e[97] * (m098 - 1))) % n;
  assign m099 = twice_mod(m098,n); assign r099 = (r098 * (1+ e[98] * (m099 - 1))) % n;
  assign m100 = twice_mod(m099,n); assign r100 = (r099 * (1+ e[99] * (m100 - 1))) % n;
  assign m101 = twice_mod(m100,n); assign r101 = (r100 * (1+ e[100] * (m101 - 1))) % n;
  assign m102 = twice_mod(m101,n); assign r102 = (r101 * (1+ e[101] * (m102 - 1))) % n;
  assign m103 = twice_mod(m102,n); assign r103 = (r102 * (1+ e[102] * (m103 - 1))) % n;
  assign m104 = twice_mod(m103,n); assign r104 = (r103 * (1+ e[103] * (m104 - 1))) % n;
  assign m105 = twice_mod(m104,n); assign r105 = (r104 * (1+ e[104] * (m105 - 1))) % n;
  assign m106 = twice_mod(m105,n); assign r106 = (r105 * (1+ e[105] * (m106 - 1))) % n;
  assign m107 = twice_mod(m106,n); assign r107 = (r106 * (1+ e[106] * (m107 - 1))) % n;
  assign m108 = twice_mod(m107,n); assign r108 = (r107 * (1+ e[107] * (m108 - 1))) % n;
  assign m109 = twice_mod(m108,n); assign r109 = (r108 * (1+ e[108] * (m109 - 1))) % n;
  assign m110 = twice_mod(m109,n); assign r110 = (r109 * (1+ e[109] * (m110 - 1))) % n;
  assign m111 = twice_mod(m110,n); assign r111 = (r110 * (1+ e[110] * (m111 - 1))) % n;
  assign m112 = twice_mod(m111,n); assign r112 = (r111 * (1+ e[111] * (m112 - 1))) % n;
  assign m113 = twice_mod(m112,n); assign r113 = (r112 * (1+ e[112] * (m113 - 1))) % n;
  assign m114 = twice_mod(m113,n); assign r114 = (r113 * (1+ e[113] * (m114 - 1))) % n;
  assign m115 = twice_mod(m114,n); assign r115 = (r114 * (1+ e[114] * (m115 - 1))) % n;
  assign m116 = twice_mod(m115,n); assign r116 = (r115 * (1+ e[115] * (m116 - 1))) % n;
  assign m117 = twice_mod(m116,n); assign r117 = (r116 * (1+ e[116] * (m117 - 1))) % n;
  assign m118 = twice_mod(m117,n); assign r118 = (r117 * (1+ e[117] * (m118 - 1))) % n;
  assign m119 = twice_mod(m118,n); assign r119 = (r118 * (1+ e[118] * (m119 - 1))) % n;
  assign m120 = twice_mod(m119,n); assign r120 = (r119 * (1+ e[119] * (m120 - 1))) % n;
  assign m121 = twice_mod(m120,n); assign r121 = (r120 * (1+ e[120] * (m121 - 1))) % n;
  assign m122 = twice_mod(m121,n); assign r122 = (r121 * (1+ e[121] * (m122 - 1))) % n;
  assign m123 = twice_mod(m122,n); assign r123 = (r122 * (1+ e[122] * (m123 - 1))) % n;
  assign m124 = twice_mod(m123,n); assign r124 = (r123 * (1+ e[123] * (m124 - 1))) % n;
  assign m125 = twice_mod(m124,n); assign r125 = (r124 * (1+ e[124] * (m125 - 1))) % n;
  assign m126 = twice_mod(m125,n); assign r126 = (r125 * (1+ e[125] * (m126 - 1))) % n;
  assign m127 = twice_mod(m126,n); assign r127 = (r126 * (1+ e[126] * (m127 - 1))) % n;
  assign m128 = twice_mod(m127,n); assign r128 = (r127 * (1+ e[127] * (m128 - 1))) % n;
  assign m129 = twice_mod(m128,n); assign r129 = (r128 * (1+ e[128] * (m129 - 1))) % n;
  assign m130 = twice_mod(m129,n); assign r130 = (r129 * (1+ e[129] * (m130 - 1))) % n;
  assign m131 = twice_mod(m130,n); assign r131 = (r130 * (1+ e[130] * (m131 - 1))) % n;
  assign m132 = twice_mod(m131,n); assign r132 = (r131 * (1+ e[131] * (m132 - 1))) % n;
  assign m133 = twice_mod(m132,n); assign r133 = (r132 * (1+ e[132] * (m133 - 1))) % n;
  assign m134 = twice_mod(m133,n); assign r134 = (r133 * (1+ e[133] * (m134 - 1))) % n;
  assign m135 = twice_mod(m134,n); assign r135 = (r134 * (1+ e[134] * (m135 - 1))) % n;
  assign m136 = twice_mod(m135,n); assign r136 = (r135 * (1+ e[135] * (m136 - 1))) % n;
  assign m137 = twice_mod(m136,n); assign r137 = (r136 * (1+ e[136] * (m137 - 1))) % n;
  assign m138 = twice_mod(m137,n); assign r138 = (r137 * (1+ e[137] * (m138 - 1))) % n;
  assign m139 = twice_mod(m138,n); assign r139 = (r138 * (1+ e[138] * (m139 - 1))) % n;
  assign m140 = twice_mod(m139,n); assign r140 = (r139 * (1+ e[139] * (m140 - 1))) % n;
  assign m141 = twice_mod(m140,n); assign r141 = (r140 * (1+ e[140] * (m141 - 1))) % n;
  assign m142 = twice_mod(m141,n); assign r142 = (r141 * (1+ e[141] * (m142 - 1))) % n;
  assign m143 = twice_mod(m142,n); assign r143 = (r142 * (1+ e[142] * (m143 - 1))) % n;
  assign m144 = twice_mod(m143,n); assign r144 = (r143 * (1+ e[143] * (m144 - 1))) % n;
  assign m145 = twice_mod(m144,n); assign r145 = (r144 * (1+ e[144] * (m145 - 1))) % n;
  assign m146 = twice_mod(m145,n); assign r146 = (r145 * (1+ e[145] * (m146 - 1))) % n;
  assign m147 = twice_mod(m146,n); assign r147 = (r146 * (1+ e[146] * (m147 - 1))) % n;
  assign m148 = twice_mod(m147,n); assign r148 = (r147 * (1+ e[147] * (m148 - 1))) % n;
  assign m149 = twice_mod(m148,n); assign r149 = (r148 * (1+ e[148] * (m149 - 1))) % n;
  assign m150 = twice_mod(m149,n); assign r150 = (r149 * (1+ e[149] * (m150 - 1))) % n;
  assign m151 = twice_mod(m150,n); assign r151 = (r150 * (1+ e[150] * (m151 - 1))) % n;
  assign m152 = twice_mod(m151,n); assign r152 = (r151 * (1+ e[151] * (m152 - 1))) % n;
  assign m153 = twice_mod(m152,n); assign r153 = (r152 * (1+ e[152] * (m153 - 1))) % n;
  assign m154 = twice_mod(m153,n); assign r154 = (r153 * (1+ e[153] * (m154 - 1))) % n;
  assign m155 = twice_mod(m154,n); assign r155 = (r154 * (1+ e[154] * (m155 - 1))) % n;
  assign m156 = twice_mod(m155,n); assign r156 = (r155 * (1+ e[155] * (m156 - 1))) % n;
  assign m157 = twice_mod(m156,n); assign r157 = (r156 * (1+ e[156] * (m157 - 1))) % n;
  assign m158 = twice_mod(m157,n); assign r158 = (r157 * (1+ e[157] * (m158 - 1))) % n;
  assign m159 = twice_mod(m158,n); assign r159 = (r158 * (1+ e[158] * (m159 - 1))) % n;
  assign m160 = twice_mod(m159,n); assign r160 = (r159 * (1+ e[159] * (m160 - 1))) % n;
  assign m161 = twice_mod(m160,n); assign r161 = (r160 * (1+ e[160] * (m161 - 1))) % n;
  assign m162 = twice_mod(m161,n); assign r162 = (r161 * (1+ e[161] * (m162 - 1))) % n;
  assign m163 = twice_mod(m162,n); assign r163 = (r162 * (1+ e[162] * (m163 - 1))) % n;
  assign m164 = twice_mod(m163,n); assign r164 = (r163 * (1+ e[163] * (m164 - 1))) % n;
  assign m165 = twice_mod(m164,n); assign r165 = (r164 * (1+ e[164] * (m165 - 1))) % n;
  assign m166 = twice_mod(m165,n); assign r166 = (r165 * (1+ e[165] * (m166 - 1))) % n;
  assign m167 = twice_mod(m166,n); assign r167 = (r166 * (1+ e[166] * (m167 - 1))) % n;
  assign m168 = twice_mod(m167,n); assign r168 = (r167 * (1+ e[167] * (m168 - 1))) % n;
  assign m169 = twice_mod(m168,n); assign r169 = (r168 * (1+ e[168] * (m169 - 1))) % n;
  assign m170 = twice_mod(m169,n); assign r170 = (r169 * (1+ e[169] * (m170 - 1))) % n;
  assign m171 = twice_mod(m170,n); assign r171 = (r170 * (1+ e[170] * (m171 - 1))) % n;
  assign m172 = twice_mod(m171,n); assign r172 = (r171 * (1+ e[171] * (m172 - 1))) % n;
  assign m173 = twice_mod(m172,n); assign r173 = (r172 * (1+ e[172] * (m173 - 1))) % n;
  assign m174 = twice_mod(m173,n); assign r174 = (r173 * (1+ e[173] * (m174 - 1))) % n;
  assign m175 = twice_mod(m174,n); assign r175 = (r174 * (1+ e[174] * (m175 - 1))) % n;
  assign m176 = twice_mod(m175,n); assign r176 = (r175 * (1+ e[175] * (m176 - 1))) % n;
  assign m177 = twice_mod(m176,n); assign r177 = (r176 * (1+ e[176] * (m177 - 1))) % n;
  assign m178 = twice_mod(m177,n); assign r178 = (r177 * (1+ e[177] * (m178 - 1))) % n;
  assign m179 = twice_mod(m178,n); assign r179 = (r178 * (1+ e[178] * (m179 - 1))) % n;
  assign m180 = twice_mod(m179,n); assign r180 = (r179 * (1+ e[179] * (m180 - 1))) % n;
  assign m181 = twice_mod(m180,n); assign r181 = (r180 * (1+ e[180] * (m181 - 1))) % n;
  assign m182 = twice_mod(m181,n); assign r182 = (r181 * (1+ e[181] * (m182 - 1))) % n;
  assign m183 = twice_mod(m182,n); assign r183 = (r182 * (1+ e[182] * (m183 - 1))) % n;
  assign m184 = twice_mod(m183,n); assign r184 = (r183 * (1+ e[183] * (m184 - 1))) % n;
  assign m185 = twice_mod(m184,n); assign r185 = (r184 * (1+ e[184] * (m185 - 1))) % n;
  assign m186 = twice_mod(m185,n); assign r186 = (r185 * (1+ e[185] * (m186 - 1))) % n;
  assign m187 = twice_mod(m186,n); assign r187 = (r186 * (1+ e[186] * (m187 - 1))) % n;
  assign m188 = twice_mod(m187,n); assign r188 = (r187 * (1+ e[187] * (m188 - 1))) % n;
  assign m189 = twice_mod(m188,n); assign r189 = (r188 * (1+ e[188] * (m189 - 1))) % n;
  assign m190 = twice_mod(m189,n); assign r190 = (r189 * (1+ e[189] * (m190 - 1))) % n;
  assign m191 = twice_mod(m190,n); assign r191 = (r190 * (1+ e[190] * (m191 - 1))) % n;
  assign m192 = twice_mod(m191,n); assign r192 = (r191 * (1+ e[191] * (m192 - 1))) % n;
  assign m193 = twice_mod(m192,n); assign r193 = (r192 * (1+ e[192] * (m193 - 1))) % n;
  assign m194 = twice_mod(m193,n); assign r194 = (r193 * (1+ e[193] * (m194 - 1))) % n;
  assign m195 = twice_mod(m194,n); assign r195 = (r194 * (1+ e[194] * (m195 - 1))) % n;
  assign m196 = twice_mod(m195,n); assign r196 = (r195 * (1+ e[195] * (m196 - 1))) % n;
  assign m197 = twice_mod(m196,n); assign r197 = (r196 * (1+ e[196] * (m197 - 1))) % n;
  assign m198 = twice_mod(m197,n); assign r198 = (r197 * (1+ e[197] * (m198 - 1))) % n;
  assign m199 = twice_mod(m198,n); assign r199 = (r198 * (1+ e[198] * (m199 - 1))) % n;
  assign m200 = twice_mod(m199,n); assign r200 = (r199 * (1+ e[199] * (m200 - 1))) % n;
  assign m201 = twice_mod(m200,n); assign r201 = (r200 * (1+ e[200] * (m201 - 1))) % n;
  assign m202 = twice_mod(m201,n); assign r202 = (r201 * (1+ e[201] * (m202 - 1))) % n;
  assign m203 = twice_mod(m202,n); assign r203 = (r202 * (1+ e[202] * (m203 - 1))) % n;
  assign m204 = twice_mod(m203,n); assign r204 = (r203 * (1+ e[203] * (m204 - 1))) % n;
  assign m205 = twice_mod(m204,n); assign r205 = (r204 * (1+ e[204] * (m205 - 1))) % n;
  assign m206 = twice_mod(m205,n); assign r206 = (r205 * (1+ e[205] * (m206 - 1))) % n;
  assign m207 = twice_mod(m206,n); assign r207 = (r206 * (1+ e[206] * (m207 - 1))) % n;
  assign m208 = twice_mod(m207,n); assign r208 = (r207 * (1+ e[207] * (m208 - 1))) % n;
  assign m209 = twice_mod(m208,n); assign r209 = (r208 * (1+ e[208] * (m209 - 1))) % n;
  assign m210 = twice_mod(m209,n); assign r210 = (r209 * (1+ e[209] * (m210 - 1))) % n;
  assign m211 = twice_mod(m210,n); assign r211 = (r210 * (1+ e[210] * (m211 - 1))) % n;
  assign m212 = twice_mod(m211,n); assign r212 = (r211 * (1+ e[211] * (m212 - 1))) % n;
  assign m213 = twice_mod(m212,n); assign r213 = (r212 * (1+ e[212] * (m213 - 1))) % n;
  assign m214 = twice_mod(m213,n); assign r214 = (r213 * (1+ e[213] * (m214 - 1))) % n;
  assign m215 = twice_mod(m214,n); assign r215 = (r214 * (1+ e[214] * (m215 - 1))) % n;
  assign m216 = twice_mod(m215,n); assign r216 = (r215 * (1+ e[215] * (m216 - 1))) % n;
  assign m217 = twice_mod(m216,n); assign r217 = (r216 * (1+ e[216] * (m217 - 1))) % n;
  assign m218 = twice_mod(m217,n); assign r218 = (r217 * (1+ e[217] * (m218 - 1))) % n;
  assign m219 = twice_mod(m218,n); assign r219 = (r218 * (1+ e[218] * (m219 - 1))) % n;
  assign m220 = twice_mod(m219,n); assign r220 = (r219 * (1+ e[219] * (m220 - 1))) % n;
  assign m221 = twice_mod(m220,n); assign r221 = (r220 * (1+ e[220] * (m221 - 1))) % n;
  assign m222 = twice_mod(m221,n); assign r222 = (r221 * (1+ e[221] * (m222 - 1))) % n;
  assign m223 = twice_mod(m222,n); assign r223 = (r222 * (1+ e[222] * (m223 - 1))) % n;
  assign m224 = twice_mod(m223,n); assign r224 = (r223 * (1+ e[223] * (m224 - 1))) % n;
  assign m225 = twice_mod(m224,n); assign r225 = (r224 * (1+ e[224] * (m225 - 1))) % n;
  assign m226 = twice_mod(m225,n); assign r226 = (r225 * (1+ e[225] * (m226 - 1))) % n;
  assign m227 = twice_mod(m226,n); assign r227 = (r226 * (1+ e[226] * (m227 - 1))) % n;
  assign m228 = twice_mod(m227,n); assign r228 = (r227 * (1+ e[227] * (m228 - 1))) % n;
  assign m229 = twice_mod(m228,n); assign r229 = (r228 * (1+ e[228] * (m229 - 1))) % n;
  assign m230 = twice_mod(m229,n); assign r230 = (r229 * (1+ e[229] * (m230 - 1))) % n;
  assign m231 = twice_mod(m230,n); assign r231 = (r230 * (1+ e[230] * (m231 - 1))) % n;
  assign m232 = twice_mod(m231,n); assign r232 = (r231 * (1+ e[231] * (m232 - 1))) % n;
  assign m233 = twice_mod(m232,n); assign r233 = (r232 * (1+ e[232] * (m233 - 1))) % n;
  assign m234 = twice_mod(m233,n); assign r234 = (r233 * (1+ e[233] * (m234 - 1))) % n;
  assign m235 = twice_mod(m234,n); assign r235 = (r234 * (1+ e[234] * (m235 - 1))) % n;
  assign m236 = twice_mod(m235,n); assign r236 = (r235 * (1+ e[235] * (m236 - 1))) % n;
  assign m237 = twice_mod(m236,n); assign r237 = (r236 * (1+ e[236] * (m237 - 1))) % n;
  assign m238 = twice_mod(m237,n); assign r238 = (r237 * (1+ e[237] * (m238 - 1))) % n;
  assign m239 = twice_mod(m238,n); assign r239 = (r238 * (1+ e[238] * (m239 - 1))) % n;
  assign m240 = twice_mod(m239,n); assign r240 = (r239 * (1+ e[239] * (m240 - 1))) % n;
  assign m241 = twice_mod(m240,n); assign r241 = (r240 * (1+ e[240] * (m241 - 1))) % n;
  assign m242 = twice_mod(m241,n); assign r242 = (r241 * (1+ e[241] * (m242 - 1))) % n;
  assign m243 = twice_mod(m242,n); assign r243 = (r242 * (1+ e[242] * (m243 - 1))) % n;
  assign m244 = twice_mod(m243,n); assign r244 = (r243 * (1+ e[243] * (m244 - 1))) % n;
  assign m245 = twice_mod(m244,n); assign r245 = (r244 * (1+ e[244] * (m245 - 1))) % n;
  assign m246 = twice_mod(m245,n); assign r246 = (r245 * (1+ e[245] * (m246 - 1))) % n;
  assign m247 = twice_mod(m246,n); assign r247 = (r246 * (1+ e[246] * (m247 - 1))) % n;
  assign m248 = twice_mod(m247,n); assign r248 = (r247 * (1+ e[247] * (m248 - 1))) % n;
  assign m249 = twice_mod(m248,n); assign r249 = (r248 * (1+ e[248] * (m249 - 1))) % n;
  assign m250 = twice_mod(m249,n); assign r250 = (r249 * (1+ e[249] * (m250 - 1))) % n;
  assign m251 = twice_mod(m250,n); assign r251 = (r250 * (1+ e[250] * (m251 - 1))) % n;
  assign m252 = twice_mod(m251,n); assign r252 = (r251 * (1+ e[251] * (m252 - 1))) % n;
  assign m253 = twice_mod(m252,n); assign r253 = (r252 * (1+ e[252] * (m253 - 1))) % n;
  assign m254 = twice_mod(m253,n); assign r254 = (r253 * (1+ e[253] * (m254 - 1))) % n;
  assign m255 = twice_mod(m254,n); assign r255 = (r254 * (1+ e[254] * (m255 - 1))) % n;
  assign m256 = twice_mod(m255,n); assign r256 = (r255 * (1+ e[255] * (m256 - 1))) % n;
  assign m257 = twice_mod(m256,n); assign r257 = (r256 * (1+ e[256] * (m257 - 1))) % n;
  assign m258 = twice_mod(m257,n); assign r258 = (r257 * (1+ e[257] * (m258 - 1))) % n;
  assign m259 = twice_mod(m258,n); assign r259 = (r258 * (1+ e[258] * (m259 - 1))) % n;
  assign m260 = twice_mod(m259,n); assign r260 = (r259 * (1+ e[259] * (m260 - 1))) % n;
  assign m261 = twice_mod(m260,n); assign r261 = (r260 * (1+ e[260] * (m261 - 1))) % n;
  assign m262 = twice_mod(m261,n); assign r262 = (r261 * (1+ e[261] * (m262 - 1))) % n;
  assign m263 = twice_mod(m262,n); assign r263 = (r262 * (1+ e[262] * (m263 - 1))) % n;
  assign m264 = twice_mod(m263,n); assign r264 = (r263 * (1+ e[263] * (m264 - 1))) % n;
  assign m265 = twice_mod(m264,n); assign r265 = (r264 * (1+ e[264] * (m265 - 1))) % n;
  assign m266 = twice_mod(m265,n); assign r266 = (r265 * (1+ e[265] * (m266 - 1))) % n;
  assign m267 = twice_mod(m266,n); assign r267 = (r266 * (1+ e[266] * (m267 - 1))) % n;
  assign m268 = twice_mod(m267,n); assign r268 = (r267 * (1+ e[267] * (m268 - 1))) % n;
  assign m269 = twice_mod(m268,n); assign r269 = (r268 * (1+ e[268] * (m269 - 1))) % n;
  assign m270 = twice_mod(m269,n); assign r270 = (r269 * (1+ e[269] * (m270 - 1))) % n;
  assign m271 = twice_mod(m270,n); assign r271 = (r270 * (1+ e[270] * (m271 - 1))) % n;
  assign m272 = twice_mod(m271,n); assign r272 = (r271 * (1+ e[271] * (m272 - 1))) % n;
  assign m273 = twice_mod(m272,n); assign r273 = (r272 * (1+ e[272] * (m273 - 1))) % n;
  assign m274 = twice_mod(m273,n); assign r274 = (r273 * (1+ e[273] * (m274 - 1))) % n;
  assign m275 = twice_mod(m274,n); assign r275 = (r274 * (1+ e[274] * (m275 - 1))) % n;
  assign m276 = twice_mod(m275,n); assign r276 = (r275 * (1+ e[275] * (m276 - 1))) % n;
  assign m277 = twice_mod(m276,n); assign r277 = (r276 * (1+ e[276] * (m277 - 1))) % n;
  assign m278 = twice_mod(m277,n); assign r278 = (r277 * (1+ e[277] * (m278 - 1))) % n;
  assign m279 = twice_mod(m278,n); assign r279 = (r278 * (1+ e[278] * (m279 - 1))) % n;
  assign m280 = twice_mod(m279,n); assign r280 = (r279 * (1+ e[279] * (m280 - 1))) % n;
  assign m281 = twice_mod(m280,n); assign r281 = (r280 * (1+ e[280] * (m281 - 1))) % n;
  assign m282 = twice_mod(m281,n); assign r282 = (r281 * (1+ e[281] * (m282 - 1))) % n;
  assign m283 = twice_mod(m282,n); assign r283 = (r282 * (1+ e[282] * (m283 - 1))) % n;
  assign m284 = twice_mod(m283,n); assign r284 = (r283 * (1+ e[283] * (m284 - 1))) % n;
  assign m285 = twice_mod(m284,n); assign r285 = (r284 * (1+ e[284] * (m285 - 1))) % n;
  assign m286 = twice_mod(m285,n); assign r286 = (r285 * (1+ e[285] * (m286 - 1))) % n;
  assign m287 = twice_mod(m286,n); assign r287 = (r286 * (1+ e[286] * (m287 - 1))) % n;
  assign m288 = twice_mod(m287,n); assign r288 = (r287 * (1+ e[287] * (m288 - 1))) % n;
  assign m289 = twice_mod(m288,n); assign r289 = (r288 * (1+ e[288] * (m289 - 1))) % n;
  assign m290 = twice_mod(m289,n); assign r290 = (r289 * (1+ e[289] * (m290 - 1))) % n;
  assign m291 = twice_mod(m290,n); assign r291 = (r290 * (1+ e[290] * (m291 - 1))) % n;
  assign m292 = twice_mod(m291,n); assign r292 = (r291 * (1+ e[291] * (m292 - 1))) % n;
  assign m293 = twice_mod(m292,n); assign r293 = (r292 * (1+ e[292] * (m293 - 1))) % n;
  assign m294 = twice_mod(m293,n); assign r294 = (r293 * (1+ e[293] * (m294 - 1))) % n;
  assign m295 = twice_mod(m294,n); assign r295 = (r294 * (1+ e[294] * (m295 - 1))) % n;
  assign m296 = twice_mod(m295,n); assign r296 = (r295 * (1+ e[295] * (m296 - 1))) % n;
  assign m297 = twice_mod(m296,n); assign r297 = (r296 * (1+ e[296] * (m297 - 1))) % n;
  assign m298 = twice_mod(m297,n); assign r298 = (r297 * (1+ e[297] * (m298 - 1))) % n;
  assign m299 = twice_mod(m298,n); assign r299 = (r298 * (1+ e[298] * (m299 - 1))) % n;
  assign m300 = twice_mod(m299,n); assign r300 = (r299 * (1+ e[299] * (m300 - 1))) % n;
  assign m301 = twice_mod(m300,n); assign r301 = (r300 * (1+ e[300] * (m301 - 1))) % n;
  assign m302 = twice_mod(m301,n); assign r302 = (r301 * (1+ e[301] * (m302 - 1))) % n;
  assign m303 = twice_mod(m302,n); assign r303 = (r302 * (1+ e[302] * (m303 - 1))) % n;
  assign m304 = twice_mod(m303,n); assign r304 = (r303 * (1+ e[303] * (m304 - 1))) % n;
  assign m305 = twice_mod(m304,n); assign r305 = (r304 * (1+ e[304] * (m305 - 1))) % n;
  assign m306 = twice_mod(m305,n); assign r306 = (r305 * (1+ e[305] * (m306 - 1))) % n;
  assign m307 = twice_mod(m306,n); assign r307 = (r306 * (1+ e[306] * (m307 - 1))) % n;
  assign m308 = twice_mod(m307,n); assign r308 = (r307 * (1+ e[307] * (m308 - 1))) % n;
  assign m309 = twice_mod(m308,n); assign r309 = (r308 * (1+ e[308] * (m309 - 1))) % n;
  assign m310 = twice_mod(m309,n); assign r310 = (r309 * (1+ e[309] * (m310 - 1))) % n;
  assign m311 = twice_mod(m310,n); assign r311 = (r310 * (1+ e[310] * (m311 - 1))) % n;
  assign m312 = twice_mod(m311,n); assign r312 = (r311 * (1+ e[311] * (m312 - 1))) % n;
  assign m313 = twice_mod(m312,n); assign r313 = (r312 * (1+ e[312] * (m313 - 1))) % n;
  assign m314 = twice_mod(m313,n); assign r314 = (r313 * (1+ e[313] * (m314 - 1))) % n;
  assign m315 = twice_mod(m314,n); assign r315 = (r314 * (1+ e[314] * (m315 - 1))) % n;
  assign m316 = twice_mod(m315,n); assign r316 = (r315 * (1+ e[315] * (m316 - 1))) % n;
  assign m317 = twice_mod(m316,n); assign r317 = (r316 * (1+ e[316] * (m317 - 1))) % n;
  assign m318 = twice_mod(m317,n); assign r318 = (r317 * (1+ e[317] * (m318 - 1))) % n;
  assign m319 = twice_mod(m318,n); assign r319 = (r318 * (1+ e[318] * (m319 - 1))) % n;
  assign m320 = twice_mod(m319,n); assign r320 = (r319 * (1+ e[319] * (m320 - 1))) % n;
  assign m321 = twice_mod(m320,n); assign r321 = (r320 * (1+ e[320] * (m321 - 1))) % n;
  assign m322 = twice_mod(m321,n); assign r322 = (r321 * (1+ e[321] * (m322 - 1))) % n;
  assign m323 = twice_mod(m322,n); assign r323 = (r322 * (1+ e[322] * (m323 - 1))) % n;
  assign m324 = twice_mod(m323,n); assign r324 = (r323 * (1+ e[323] * (m324 - 1))) % n;
  assign m325 = twice_mod(m324,n); assign r325 = (r324 * (1+ e[324] * (m325 - 1))) % n;
  assign m326 = twice_mod(m325,n); assign r326 = (r325 * (1+ e[325] * (m326 - 1))) % n;
  assign m327 = twice_mod(m326,n); assign r327 = (r326 * (1+ e[326] * (m327 - 1))) % n;
  assign m328 = twice_mod(m327,n); assign r328 = (r327 * (1+ e[327] * (m328 - 1))) % n;
  assign m329 = twice_mod(m328,n); assign r329 = (r328 * (1+ e[328] * (m329 - 1))) % n;
  assign m330 = twice_mod(m329,n); assign r330 = (r329 * (1+ e[329] * (m330 - 1))) % n;
  assign m331 = twice_mod(m330,n); assign r331 = (r330 * (1+ e[330] * (m331 - 1))) % n;
  assign m332 = twice_mod(m331,n); assign r332 = (r331 * (1+ e[331] * (m332 - 1))) % n;
  assign m333 = twice_mod(m332,n); assign r333 = (r332 * (1+ e[332] * (m333 - 1))) % n;
  assign m334 = twice_mod(m333,n); assign r334 = (r333 * (1+ e[333] * (m334 - 1))) % n;
  assign m335 = twice_mod(m334,n); assign r335 = (r334 * (1+ e[334] * (m335 - 1))) % n;
  assign m336 = twice_mod(m335,n); assign r336 = (r335 * (1+ e[335] * (m336 - 1))) % n;
  assign m337 = twice_mod(m336,n); assign r337 = (r336 * (1+ e[336] * (m337 - 1))) % n;
  assign m338 = twice_mod(m337,n); assign r338 = (r337 * (1+ e[337] * (m338 - 1))) % n;
  assign m339 = twice_mod(m338,n); assign r339 = (r338 * (1+ e[338] * (m339 - 1))) % n;
  assign m340 = twice_mod(m339,n); assign r340 = (r339 * (1+ e[339] * (m340 - 1))) % n;
  assign m341 = twice_mod(m340,n); assign r341 = (r340 * (1+ e[340] * (m341 - 1))) % n;
  assign m342 = twice_mod(m341,n); assign r342 = (r341 * (1+ e[341] * (m342 - 1))) % n;
  assign m343 = twice_mod(m342,n); assign r343 = (r342 * (1+ e[342] * (m343 - 1))) % n;
  assign m344 = twice_mod(m343,n); assign r344 = (r343 * (1+ e[343] * (m344 - 1))) % n;
  assign m345 = twice_mod(m344,n); assign r345 = (r344 * (1+ e[344] * (m345 - 1))) % n;
  assign m346 = twice_mod(m345,n); assign r346 = (r345 * (1+ e[345] * (m346 - 1))) % n;
  assign m347 = twice_mod(m346,n); assign r347 = (r346 * (1+ e[346] * (m347 - 1))) % n;
  assign m348 = twice_mod(m347,n); assign r348 = (r347 * (1+ e[347] * (m348 - 1))) % n;
  assign m349 = twice_mod(m348,n); assign r349 = (r348 * (1+ e[348] * (m349 - 1))) % n;
  assign m350 = twice_mod(m349,n); assign r350 = (r349 * (1+ e[349] * (m350 - 1))) % n;
  assign m351 = twice_mod(m350,n); assign r351 = (r350 * (1+ e[350] * (m351 - 1))) % n;
  assign m352 = twice_mod(m351,n); assign r352 = (r351 * (1+ e[351] * (m352 - 1))) % n;
  assign m353 = twice_mod(m352,n); assign r353 = (r352 * (1+ e[352] * (m353 - 1))) % n;
  assign m354 = twice_mod(m353,n); assign r354 = (r353 * (1+ e[353] * (m354 - 1))) % n;
  assign m355 = twice_mod(m354,n); assign r355 = (r354 * (1+ e[354] * (m355 - 1))) % n;
  assign m356 = twice_mod(m355,n); assign r356 = (r355 * (1+ e[355] * (m356 - 1))) % n;
  assign m357 = twice_mod(m356,n); assign r357 = (r356 * (1+ e[356] * (m357 - 1))) % n;
  assign m358 = twice_mod(m357,n); assign r358 = (r357 * (1+ e[357] * (m358 - 1))) % n;
  assign m359 = twice_mod(m358,n); assign r359 = (r358 * (1+ e[358] * (m359 - 1))) % n;
  assign m360 = twice_mod(m359,n); assign r360 = (r359 * (1+ e[359] * (m360 - 1))) % n;
  assign m361 = twice_mod(m360,n); assign r361 = (r360 * (1+ e[360] * (m361 - 1))) % n;
  assign m362 = twice_mod(m361,n); assign r362 = (r361 * (1+ e[361] * (m362 - 1))) % n;
  assign m363 = twice_mod(m362,n); assign r363 = (r362 * (1+ e[362] * (m363 - 1))) % n;
  assign m364 = twice_mod(m363,n); assign r364 = (r363 * (1+ e[363] * (m364 - 1))) % n;
  assign m365 = twice_mod(m364,n); assign r365 = (r364 * (1+ e[364] * (m365 - 1))) % n;
  assign m366 = twice_mod(m365,n); assign r366 = (r365 * (1+ e[365] * (m366 - 1))) % n;
  assign m367 = twice_mod(m366,n); assign r367 = (r366 * (1+ e[366] * (m367 - 1))) % n;
  assign m368 = twice_mod(m367,n); assign r368 = (r367 * (1+ e[367] * (m368 - 1))) % n;
  assign m369 = twice_mod(m368,n); assign r369 = (r368 * (1+ e[368] * (m369 - 1))) % n;
  assign m370 = twice_mod(m369,n); assign r370 = (r369 * (1+ e[369] * (m370 - 1))) % n;
  assign m371 = twice_mod(m370,n); assign r371 = (r370 * (1+ e[370] * (m371 - 1))) % n;
  assign m372 = twice_mod(m371,n); assign r372 = (r371 * (1+ e[371] * (m372 - 1))) % n;
  assign m373 = twice_mod(m372,n); assign r373 = (r372 * (1+ e[372] * (m373 - 1))) % n;
  assign m374 = twice_mod(m373,n); assign r374 = (r373 * (1+ e[373] * (m374 - 1))) % n;
  assign m375 = twice_mod(m374,n); assign r375 = (r374 * (1+ e[374] * (m375 - 1))) % n;
  assign m376 = twice_mod(m375,n); assign r376 = (r375 * (1+ e[375] * (m376 - 1))) % n;
  assign m377 = twice_mod(m376,n); assign r377 = (r376 * (1+ e[376] * (m377 - 1))) % n;
  assign m378 = twice_mod(m377,n); assign r378 = (r377 * (1+ e[377] * (m378 - 1))) % n;
  assign m379 = twice_mod(m378,n); assign r379 = (r378 * (1+ e[378] * (m379 - 1))) % n;
  assign m380 = twice_mod(m379,n); assign r380 = (r379 * (1+ e[379] * (m380 - 1))) % n;
  assign m381 = twice_mod(m380,n); assign r381 = (r380 * (1+ e[380] * (m381 - 1))) % n;
  assign m382 = twice_mod(m381,n); assign r382 = (r381 * (1+ e[381] * (m382 - 1))) % n;
  assign m383 = twice_mod(m382,n); assign r383 = (r382 * (1+ e[382] * (m383 - 1))) % n;
  assign m384 = twice_mod(m383,n); assign r384 = (r383 * (1+ e[383] * (m384 - 1))) % n;
  assign m385 = twice_mod(m384,n); assign r385 = (r384 * (1+ e[384] * (m385 - 1))) % n;
  assign m386 = twice_mod(m385,n); assign r386 = (r385 * (1+ e[385] * (m386 - 1))) % n;
  assign m387 = twice_mod(m386,n); assign r387 = (r386 * (1+ e[386] * (m387 - 1))) % n;
  assign m388 = twice_mod(m387,n); assign r388 = (r387 * (1+ e[387] * (m388 - 1))) % n;
  assign m389 = twice_mod(m388,n); assign r389 = (r388 * (1+ e[388] * (m389 - 1))) % n;
  assign m390 = twice_mod(m389,n); assign r390 = (r389 * (1+ e[389] * (m390 - 1))) % n;
  assign m391 = twice_mod(m390,n); assign r391 = (r390 * (1+ e[390] * (m391 - 1))) % n;
  assign m392 = twice_mod(m391,n); assign r392 = (r391 * (1+ e[391] * (m392 - 1))) % n;
  assign m393 = twice_mod(m392,n); assign r393 = (r392 * (1+ e[392] * (m393 - 1))) % n;
  assign m394 = twice_mod(m393,n); assign r394 = (r393 * (1+ e[393] * (m394 - 1))) % n;
  assign m395 = twice_mod(m394,n); assign r395 = (r394 * (1+ e[394] * (m395 - 1))) % n;
  assign m396 = twice_mod(m395,n); assign r396 = (r395 * (1+ e[395] * (m396 - 1))) % n;
  assign m397 = twice_mod(m396,n); assign r397 = (r396 * (1+ e[396] * (m397 - 1))) % n;
  assign m398 = twice_mod(m397,n); assign r398 = (r397 * (1+ e[397] * (m398 - 1))) % n;
  assign m399 = twice_mod(m398,n); assign r399 = (r398 * (1+ e[398] * (m399 - 1))) % n;
  assign m400 = twice_mod(m399,n); assign r400 = (r399 * (1+ e[399] * (m400 - 1))) % n;
  assign m401 = twice_mod(m400,n); assign r401 = (r400 * (1+ e[400] * (m401 - 1))) % n;
  assign m402 = twice_mod(m401,n); assign r402 = (r401 * (1+ e[401] * (m402 - 1))) % n;
  assign m403 = twice_mod(m402,n); assign r403 = (r402 * (1+ e[402] * (m403 - 1))) % n;
  assign m404 = twice_mod(m403,n); assign r404 = (r403 * (1+ e[403] * (m404 - 1))) % n;
  assign m405 = twice_mod(m404,n); assign r405 = (r404 * (1+ e[404] * (m405 - 1))) % n;
  assign m406 = twice_mod(m405,n); assign r406 = (r405 * (1+ e[405] * (m406 - 1))) % n;
  assign m407 = twice_mod(m406,n); assign r407 = (r406 * (1+ e[406] * (m407 - 1))) % n;
  assign m408 = twice_mod(m407,n); assign r408 = (r407 * (1+ e[407] * (m408 - 1))) % n;
  assign m409 = twice_mod(m408,n); assign r409 = (r408 * (1+ e[408] * (m409 - 1))) % n;
  assign m410 = twice_mod(m409,n); assign r410 = (r409 * (1+ e[409] * (m410 - 1))) % n;
  assign m411 = twice_mod(m410,n); assign r411 = (r410 * (1+ e[410] * (m411 - 1))) % n;
  assign m412 = twice_mod(m411,n); assign r412 = (r411 * (1+ e[411] * (m412 - 1))) % n;
  assign m413 = twice_mod(m412,n); assign r413 = (r412 * (1+ e[412] * (m413 - 1))) % n;
  assign m414 = twice_mod(m413,n); assign r414 = (r413 * (1+ e[413] * (m414 - 1))) % n;
  assign m415 = twice_mod(m414,n); assign r415 = (r414 * (1+ e[414] * (m415 - 1))) % n;
  assign m416 = twice_mod(m415,n); assign r416 = (r415 * (1+ e[415] * (m416 - 1))) % n;
  assign m417 = twice_mod(m416,n); assign r417 = (r416 * (1+ e[416] * (m417 - 1))) % n;
  assign m418 = twice_mod(m417,n); assign r418 = (r417 * (1+ e[417] * (m418 - 1))) % n;
  assign m419 = twice_mod(m418,n); assign r419 = (r418 * (1+ e[418] * (m419 - 1))) % n;
  assign m420 = twice_mod(m419,n); assign r420 = (r419 * (1+ e[419] * (m420 - 1))) % n;
  assign m421 = twice_mod(m420,n); assign r421 = (r420 * (1+ e[420] * (m421 - 1))) % n;
  assign m422 = twice_mod(m421,n); assign r422 = (r421 * (1+ e[421] * (m422 - 1))) % n;
  assign m423 = twice_mod(m422,n); assign r423 = (r422 * (1+ e[422] * (m423 - 1))) % n;
  assign m424 = twice_mod(m423,n); assign r424 = (r423 * (1+ e[423] * (m424 - 1))) % n;
  assign m425 = twice_mod(m424,n); assign r425 = (r424 * (1+ e[424] * (m425 - 1))) % n;
  assign m426 = twice_mod(m425,n); assign r426 = (r425 * (1+ e[425] * (m426 - 1))) % n;
  assign m427 = twice_mod(m426,n); assign r427 = (r426 * (1+ e[426] * (m427 - 1))) % n;
  assign m428 = twice_mod(m427,n); assign r428 = (r427 * (1+ e[427] * (m428 - 1))) % n;
  assign m429 = twice_mod(m428,n); assign r429 = (r428 * (1+ e[428] * (m429 - 1))) % n;
  assign m430 = twice_mod(m429,n); assign r430 = (r429 * (1+ e[429] * (m430 - 1))) % n;
  assign m431 = twice_mod(m430,n); assign r431 = (r430 * (1+ e[430] * (m431 - 1))) % n;
  assign m432 = twice_mod(m431,n); assign r432 = (r431 * (1+ e[431] * (m432 - 1))) % n;
  assign m433 = twice_mod(m432,n); assign r433 = (r432 * (1+ e[432] * (m433 - 1))) % n;
  assign m434 = twice_mod(m433,n); assign r434 = (r433 * (1+ e[433] * (m434 - 1))) % n;
  assign m435 = twice_mod(m434,n); assign r435 = (r434 * (1+ e[434] * (m435 - 1))) % n;
  assign m436 = twice_mod(m435,n); assign r436 = (r435 * (1+ e[435] * (m436 - 1))) % n;
  assign m437 = twice_mod(m436,n); assign r437 = (r436 * (1+ e[436] * (m437 - 1))) % n;
  assign m438 = twice_mod(m437,n); assign r438 = (r437 * (1+ e[437] * (m438 - 1))) % n;
  assign m439 = twice_mod(m438,n); assign r439 = (r438 * (1+ e[438] * (m439 - 1))) % n;
  assign m440 = twice_mod(m439,n); assign r440 = (r439 * (1+ e[439] * (m440 - 1))) % n;
  assign m441 = twice_mod(m440,n); assign r441 = (r440 * (1+ e[440] * (m441 - 1))) % n;
  assign m442 = twice_mod(m441,n); assign r442 = (r441 * (1+ e[441] * (m442 - 1))) % n;
  assign m443 = twice_mod(m442,n); assign r443 = (r442 * (1+ e[442] * (m443 - 1))) % n;
  assign m444 = twice_mod(m443,n); assign r444 = (r443 * (1+ e[443] * (m444 - 1))) % n;
  assign m445 = twice_mod(m444,n); assign r445 = (r444 * (1+ e[444] * (m445 - 1))) % n;
  assign m446 = twice_mod(m445,n); assign r446 = (r445 * (1+ e[445] * (m446 - 1))) % n;
  assign m447 = twice_mod(m446,n); assign r447 = (r446 * (1+ e[446] * (m447 - 1))) % n;
  assign m448 = twice_mod(m447,n); assign r448 = (r447 * (1+ e[447] * (m448 - 1))) % n;
  assign m449 = twice_mod(m448,n); assign r449 = (r448 * (1+ e[448] * (m449 - 1))) % n;
  assign m450 = twice_mod(m449,n); assign r450 = (r449 * (1+ e[449] * (m450 - 1))) % n;
  assign m451 = twice_mod(m450,n); assign r451 = (r450 * (1+ e[450] * (m451 - 1))) % n;
  assign m452 = twice_mod(m451,n); assign r452 = (r451 * (1+ e[451] * (m452 - 1))) % n;
  assign m453 = twice_mod(m452,n); assign r453 = (r452 * (1+ e[452] * (m453 - 1))) % n;
  assign m454 = twice_mod(m453,n); assign r454 = (r453 * (1+ e[453] * (m454 - 1))) % n;
  assign m455 = twice_mod(m454,n); assign r455 = (r454 * (1+ e[454] * (m455 - 1))) % n;
  assign m456 = twice_mod(m455,n); assign r456 = (r455 * (1+ e[455] * (m456 - 1))) % n;
  assign m457 = twice_mod(m456,n); assign r457 = (r456 * (1+ e[456] * (m457 - 1))) % n;
  assign m458 = twice_mod(m457,n); assign r458 = (r457 * (1+ e[457] * (m458 - 1))) % n;
  assign m459 = twice_mod(m458,n); assign r459 = (r458 * (1+ e[458] * (m459 - 1))) % n;
  assign m460 = twice_mod(m459,n); assign r460 = (r459 * (1+ e[459] * (m460 - 1))) % n;
  assign m461 = twice_mod(m460,n); assign r461 = (r460 * (1+ e[460] * (m461 - 1))) % n;
  assign m462 = twice_mod(m461,n); assign r462 = (r461 * (1+ e[461] * (m462 - 1))) % n;
  assign m463 = twice_mod(m462,n); assign r463 = (r462 * (1+ e[462] * (m463 - 1))) % n;
  assign m464 = twice_mod(m463,n); assign r464 = (r463 * (1+ e[463] * (m464 - 1))) % n;
  assign m465 = twice_mod(m464,n); assign r465 = (r464 * (1+ e[464] * (m465 - 1))) % n;
  assign m466 = twice_mod(m465,n); assign r466 = (r465 * (1+ e[465] * (m466 - 1))) % n;
  assign m467 = twice_mod(m466,n); assign r467 = (r466 * (1+ e[466] * (m467 - 1))) % n;
  assign m468 = twice_mod(m467,n); assign r468 = (r467 * (1+ e[467] * (m468 - 1))) % n;
  assign m469 = twice_mod(m468,n); assign r469 = (r468 * (1+ e[468] * (m469 - 1))) % n;
  assign m470 = twice_mod(m469,n); assign r470 = (r469 * (1+ e[469] * (m470 - 1))) % n;
  assign m471 = twice_mod(m470,n); assign r471 = (r470 * (1+ e[470] * (m471 - 1))) % n;
  assign m472 = twice_mod(m471,n); assign r472 = (r471 * (1+ e[471] * (m472 - 1))) % n;
  assign m473 = twice_mod(m472,n); assign r473 = (r472 * (1+ e[472] * (m473 - 1))) % n;
  assign m474 = twice_mod(m473,n); assign r474 = (r473 * (1+ e[473] * (m474 - 1))) % n;
  assign m475 = twice_mod(m474,n); assign r475 = (r474 * (1+ e[474] * (m475 - 1))) % n;
  assign m476 = twice_mod(m475,n); assign r476 = (r475 * (1+ e[475] * (m476 - 1))) % n;
  assign m477 = twice_mod(m476,n); assign r477 = (r476 * (1+ e[476] * (m477 - 1))) % n;
  assign m478 = twice_mod(m477,n); assign r478 = (r477 * (1+ e[477] * (m478 - 1))) % n;
  assign m479 = twice_mod(m478,n); assign r479 = (r478 * (1+ e[478] * (m479 - 1))) % n;
  assign m480 = twice_mod(m479,n); assign r480 = (r479 * (1+ e[479] * (m480 - 1))) % n;
  assign m481 = twice_mod(m480,n); assign r481 = (r480 * (1+ e[480] * (m481 - 1))) % n;
  assign m482 = twice_mod(m481,n); assign r482 = (r481 * (1+ e[481] * (m482 - 1))) % n;
  assign m483 = twice_mod(m482,n); assign r483 = (r482 * (1+ e[482] * (m483 - 1))) % n;
  assign m484 = twice_mod(m483,n); assign r484 = (r483 * (1+ e[483] * (m484 - 1))) % n;
  assign m485 = twice_mod(m484,n); assign r485 = (r484 * (1+ e[484] * (m485 - 1))) % n;
  assign m486 = twice_mod(m485,n); assign r486 = (r485 * (1+ e[485] * (m486 - 1))) % n;
  assign m487 = twice_mod(m486,n); assign r487 = (r486 * (1+ e[486] * (m487 - 1))) % n;
  assign m488 = twice_mod(m487,n); assign r488 = (r487 * (1+ e[487] * (m488 - 1))) % n;
  assign m489 = twice_mod(m488,n); assign r489 = (r488 * (1+ e[488] * (m489 - 1))) % n;
  assign m490 = twice_mod(m489,n); assign r490 = (r489 * (1+ e[489] * (m490 - 1))) % n;
  assign m491 = twice_mod(m490,n); assign r491 = (r490 * (1+ e[490] * (m491 - 1))) % n;
  assign m492 = twice_mod(m491,n); assign r492 = (r491 * (1+ e[491] * (m492 - 1))) % n;
  assign m493 = twice_mod(m492,n); assign r493 = (r492 * (1+ e[492] * (m493 - 1))) % n;
  assign m494 = twice_mod(m493,n); assign r494 = (r493 * (1+ e[493] * (m494 - 1))) % n;
  assign m495 = twice_mod(m494,n); assign r495 = (r494 * (1+ e[494] * (m495 - 1))) % n;
  assign m496 = twice_mod(m495,n); assign r496 = (r495 * (1+ e[495] * (m496 - 1))) % n;
  assign m497 = twice_mod(m496,n); assign r497 = (r496 * (1+ e[496] * (m497 - 1))) % n;
  assign m498 = twice_mod(m497,n); assign r498 = (r497 * (1+ e[497] * (m498 - 1))) % n;
  assign m499 = twice_mod(m498,n); assign r499 = (r498 * (1+ e[498] * (m499 - 1))) % n;
  assign m500 = twice_mod(m499,n); assign r500 = (r499 * (1+ e[499] * (m500 - 1))) % n;
  assign m501 = twice_mod(m500,n); assign r501 = (r500 * (1+ e[500] * (m501 - 1))) % n;
  assign m502 = twice_mod(m501,n); assign r502 = (r501 * (1+ e[501] * (m502 - 1))) % n;
  assign m503 = twice_mod(m502,n); assign r503 = (r502 * (1+ e[502] * (m503 - 1))) % n;
  assign m504 = twice_mod(m503,n); assign r504 = (r503 * (1+ e[503] * (m504 - 1))) % n;
  assign m505 = twice_mod(m504,n); assign r505 = (r504 * (1+ e[504] * (m505 - 1))) % n;
  assign m506 = twice_mod(m505,n); assign r506 = (r505 * (1+ e[505] * (m506 - 1))) % n;
  assign m507 = twice_mod(m506,n); assign r507 = (r506 * (1+ e[506] * (m507 - 1))) % n;
  assign m508 = twice_mod(m507,n); assign r508 = (r507 * (1+ e[507] * (m508 - 1))) % n;
  assign m509 = twice_mod(m508,n); assign r509 = (r508 * (1+ e[508] * (m509 - 1))) % n;
  assign m510 = twice_mod(m509,n); assign r510 = (r509 * (1+ e[509] * (m510 - 1))) % n;
  assign m511 = twice_mod(m510,n); assign r511 = (r510 * (1+ e[510] * (m511 - 1))) % n;
  assign m512 = twice_mod(m511,n); assign r512 = (r511 * (1+ e[511] * (m512 - 1))) % n;

  assign r = r512;

  function [511:0] twice_mod;
    input [511:0] m, n;
    twice_mod = (m * m) % n;
  endfunction

endmodule





module test;
  reg  [0:511]e,n,m;
  wire [0:511]r;

  initial begin
    #10
      n  <= 512'hdeadbeefdeadbeefdeadbeefdeadbeefdeadbeefdeadbeefdeadbeefdeadbeef;
      m  <= 512'hd000000000000000000000000000000000000000000000000000000000000001;
//      n  <= 16;
//      m  <= 3;
      e  <= 3;
    #1000 e <= 4;
  end

  modexp1 aab(e,n,m,r);

  initial begin
    $monitor ($stime , " hello world e:%h n:%h m:%h r:%h ",e,n,m,r);
//    $monitor ($stime , " hello world aab.e:%h aab.n:%h aab.m:%h aab.r:%h ",aab.e,aab.n,aab.m,aab.r);
    $monitor ($stime , " r001 %h r002 %h r003 %h",aab.r001,aab.r002,aab.r003);
//    $monitor ($stime , " m001 %h m002 %h m003 %h",aab.m001,aab.m002,aab.m003);
//    $monitor ($stime , " e[1] %h e[2] %h e[3] %h",aab.e[0],aab.e[1],aab.e[2]);
  end

endmodule


